magic
tech sky130A
magscale 1 2
timestamp 1624402156
<< nwell >>
rect 14730 660108 64962 661110
rect 14730 660034 64841 660108
rect 82888 660083 133067 660649
rect 83408 660052 119178 660083
rect 14730 659150 14782 660034
rect 28401 659941 28758 659982
rect 83408 659846 112858 660052
rect 124441 660015 133067 660083
<< pwell >>
rect 371257 636863 371689 637515
<< nsubdiff >>
rect 14777 660157 14801 660354
rect 21672 660157 21696 660354
rect 23064 660169 23088 660375
rect 28678 660169 28702 660375
rect 28954 660172 28978 660367
rect 34940 660172 34964 660367
rect 35514 660153 35538 660369
rect 63779 660153 63803 660369
rect 84063 660216 84087 660457
rect 112239 660216 112263 660457
rect 112659 660076 112683 660241
rect 119084 660076 119108 660241
rect 119365 660188 119389 660416
rect 124370 660188 124394 660416
rect 124754 660180 124778 660424
rect 132540 660180 132564 660424
<< nsubdiffcont >>
rect 14801 660157 21672 660354
rect 23088 660169 28678 660375
rect 28978 660172 34940 660367
rect 35538 660153 63779 660369
rect 84087 660216 112239 660457
rect 112683 660076 119084 660241
rect 119389 660188 124370 660416
rect 124778 660180 132540 660424
<< locali >>
rect 14785 660157 14801 660354
rect 21672 660157 21688 660354
rect 23072 660169 23088 660375
rect 28678 660169 28694 660375
rect 28962 660172 28978 660367
rect 34940 660172 34956 660367
rect 35522 660153 35538 660369
rect 63779 660153 63795 660369
rect 84071 660216 84087 660457
rect 112239 660216 112255 660457
rect 112667 660076 112683 660241
rect 119084 660076 119100 660241
rect 119373 660188 119389 660416
rect 124370 660188 124386 660416
<< viali >>
rect 14801 660157 21672 660354
rect 23088 660169 28678 660375
rect 28978 660172 34940 660367
rect 35538 660153 63779 660369
rect 84087 660216 112239 660457
rect 112683 660076 119084 660241
rect 119389 660188 124370 660416
rect 124762 660180 124778 660424
rect 124778 660180 132540 660424
rect 132540 660180 132556 660424
<< metal1 >>
rect 202956 687835 202966 688225
rect 206549 687835 206559 688225
rect 207113 687795 207123 688222
rect 210595 687795 210605 688222
rect 211166 687819 211176 688246
rect 214648 687819 214658 688246
rect 223050 688060 223060 688186
rect 223016 687894 223060 688060
rect 223050 687834 223060 687894
rect 226864 688060 226874 688186
rect 226864 687894 226915 688060
rect 226864 687834 226874 687894
rect 227267 687846 227277 688273
rect 230749 687846 230759 688273
rect 231320 687855 231330 688282
rect 234802 687855 234812 688282
rect 235302 687865 235312 688292
rect 238784 687865 238794 688292
rect 239323 687860 239333 688287
rect 242805 687860 242815 688287
rect 243362 687858 243372 688285
rect 246844 687858 246854 688285
rect 202763 685044 202773 685354
rect 247145 685044 247155 685354
rect 83775 660472 112339 660489
rect 23004 660431 64063 660453
rect 23004 660397 23042 660431
rect 21700 660392 23042 660397
rect 14751 660388 23042 660392
rect 14751 660354 14834 660388
rect 14751 660157 14801 660354
rect 14751 660121 14834 660157
rect 14751 660101 23042 660121
rect 64025 660101 64063 660431
rect 14751 660070 64063 660101
rect 14751 660012 21718 660070
rect 23004 660030 64063 660070
rect 23037 660018 28912 660030
rect 14751 659692 14783 660012
rect 83746 659999 83756 660472
rect 112324 660409 112339 660472
rect 119184 660445 133061 660493
rect 119184 660416 120252 660445
rect 112324 660408 112754 660409
rect 119106 660408 119389 660416
rect 112324 660332 119389 660408
rect 112324 660010 112657 660332
rect 119074 660241 119389 660332
rect 119084 660188 119389 660241
rect 119084 660106 120252 660188
rect 133038 660416 133061 660445
rect 133038 660106 133067 660416
rect 119084 660076 133067 660106
rect 112324 659999 112334 660010
rect 112601 659953 112657 660010
rect 119074 660062 133067 660076
rect 119074 659953 119177 660062
rect 125643 660015 133067 660062
rect 112601 659944 119177 659953
rect 157073 659472 157083 659901
rect 198006 659472 198016 659901
rect 12990 659376 14703 659415
rect 12990 659103 13065 659376
rect 14624 659270 14703 659376
rect 133071 659270 133081 659303
rect 14624 659204 14991 659270
rect 132917 659204 133081 659270
rect 14624 659103 14703 659204
rect 133071 659175 133081 659204
rect 133354 659175 133364 659303
rect 12990 659070 14703 659103
rect 66160 658984 66170 659137
rect 64423 658604 66170 658984
rect 63068 658320 66170 658604
rect 64423 657999 66170 658320
rect 66160 657870 66170 657999
rect 68582 658984 68592 659137
rect 68582 657999 68603 658984
rect 79846 658972 83253 658973
rect 68582 657870 68592 657999
rect 79838 657985 79848 658972
rect 82308 658604 83253 658972
rect 206575 658728 206585 658758
rect 206248 658662 206585 658728
rect 206575 658630 206585 658662
rect 206858 658630 206868 658758
rect 82308 658320 84035 658604
rect 149997 658524 156268 658555
rect 82308 657988 83253 658320
rect 82308 657985 82318 657988
rect 21150 657532 21160 657665
rect 23640 657532 23650 657665
rect 64013 657266 64962 657593
rect 34969 657163 34979 657242
rect 35060 657163 35070 657242
rect 34989 656786 35045 657163
rect 34964 656680 34974 656786
rect 35066 656680 35076 656786
rect 64135 656771 64962 657266
rect 64163 656761 64962 656771
rect 64457 656747 64962 656761
rect 82894 657275 83827 657583
rect 124326 657529 124336 657669
rect 126700 657529 126710 657669
rect 149987 657395 149997 658524
rect 152333 658062 156268 658524
rect 152333 657778 157347 658062
rect 152333 657395 156268 657778
rect 149997 657379 156268 657395
rect 82894 656573 83702 657275
rect 112660 657160 112670 657243
rect 112802 657160 112812 657243
rect 112685 656533 112741 657160
rect 156207 656708 157418 657036
rect 197704 657001 197714 657125
rect 199942 657001 199952 657125
rect 112626 656348 112636 656533
rect 112797 656348 112807 656533
rect 156207 656248 156786 656708
rect 186130 656623 186140 656702
rect 186225 656623 186235 656702
rect 186152 656414 186208 656623
rect 186119 656316 186129 656414
rect 186241 656316 186251 656414
rect 12125 655528 13406 655533
rect 12125 655200 14468 655528
rect 133382 655200 135242 655528
rect 12125 652870 13406 655200
rect 134093 653281 135239 655200
rect 207475 654986 208245 655013
rect 206694 654658 208245 654986
rect 12125 651670 15784 652870
rect 132088 652146 135239 653281
rect 207475 652403 208245 654658
rect 132558 652135 135239 652146
rect 12125 651669 15583 651670
rect 12125 651650 13406 651669
rect 205405 651403 208245 652403
rect 205405 651383 207885 651403
rect 124847 637057 124857 637281
rect 125442 637057 125452 637281
<< via1 >>
rect 202966 687835 206549 688225
rect 207123 687795 210595 688222
rect 211176 687819 214648 688246
rect 223060 687834 226864 688186
rect 227277 687846 230749 688273
rect 231330 687855 234802 688282
rect 235312 687865 238784 688292
rect 239333 687860 242805 688287
rect 243372 687858 246844 688285
rect 202773 685044 247145 685354
rect 23042 660388 64025 660431
rect 14834 660375 64025 660388
rect 14834 660354 23088 660375
rect 14834 660157 21672 660354
rect 21672 660169 23088 660354
rect 23088 660169 28678 660375
rect 28678 660369 64025 660375
rect 28678 660367 35538 660369
rect 28678 660172 28978 660367
rect 28978 660172 34940 660367
rect 34940 660172 35538 660367
rect 28678 660169 35538 660172
rect 21672 660157 35538 660169
rect 14834 660153 35538 660157
rect 35538 660153 63779 660369
rect 63779 660153 64025 660369
rect 14834 660121 64025 660153
rect 23042 660101 64025 660121
rect 83756 660457 112324 660472
rect 83756 660216 84087 660457
rect 84087 660216 112239 660457
rect 112239 660216 112324 660457
rect 120252 660424 133038 660445
rect 120252 660416 124762 660424
rect 83756 659999 112324 660216
rect 112657 660241 119074 660332
rect 112657 660076 112683 660241
rect 112683 660076 119074 660241
rect 120252 660188 124370 660416
rect 124370 660188 124762 660416
rect 120252 660180 124762 660188
rect 124762 660180 132556 660424
rect 132556 660180 133038 660424
rect 120252 660106 133038 660180
rect 112657 659953 119074 660076
rect 157083 659472 198006 659901
rect 13065 659103 14624 659376
rect 133081 659175 133354 659303
rect 66170 657870 68582 659137
rect 79848 657985 82308 658972
rect 206585 658630 206858 658758
rect 21160 657532 23640 657665
rect 34979 657163 35060 657242
rect 34974 656680 35066 656786
rect 124336 657529 126700 657669
rect 149997 657395 152333 658524
rect 112670 657160 112802 657243
rect 197714 657001 199942 657125
rect 112636 656348 112797 656533
rect 186140 656623 186225 656702
rect 186129 656316 186241 656414
rect 124857 637057 125442 637281
<< metal2 >>
rect 211169 688703 214642 688713
rect 207123 688623 210596 688633
rect 198295 688226 199269 688229
rect 202966 688226 206549 688235
rect 198295 688225 206549 688226
rect 198295 688219 202966 688225
rect 199269 687835 202966 688219
rect 199269 687830 206549 687835
rect 198295 687825 206549 687830
rect 198295 687820 199269 687825
rect 235312 688693 238785 688703
rect 231330 688683 234803 688693
rect 227277 688664 230750 688674
rect 214642 688246 214648 688256
rect 211169 687865 211176 687875
rect 223060 688186 226864 688196
rect 223060 687824 226864 687834
rect 235312 687855 238785 687865
rect 239333 688688 242806 688698
rect 231330 687845 234803 687855
rect 239333 687850 242806 687860
rect 243372 688686 246845 688696
rect 243372 687848 246845 687858
rect 227277 687826 230750 687836
rect 211176 687809 214648 687819
rect 207123 687785 210596 687795
rect 202773 685354 247145 685364
rect 202773 685034 202780 685044
rect 247142 685034 247145 685044
rect 202780 684701 247142 684711
rect 83765 660846 124085 660856
rect 23042 660657 64025 660667
rect 14834 660388 23042 660398
rect 14834 660111 23042 660121
rect 23042 660091 64025 660101
rect 83756 660472 83765 660482
rect 157083 660502 197708 660512
rect 124085 660445 133038 660455
rect 112324 659999 112657 660179
rect 83756 659989 112324 659999
rect 119074 660106 120252 660179
rect 119074 660096 133038 660106
rect 119074 659999 120418 660096
rect 112657 659943 119074 659953
rect 197708 659901 198006 659911
rect 2509 659760 14155 659826
rect 2509 658727 2671 659760
rect 5073 659386 14155 659760
rect 133210 659558 140004 659630
rect 5073 659376 14624 659386
rect 5073 659103 13065 659376
rect 133210 659313 137580 659558
rect 133081 659303 137580 659313
rect 133354 659175 137580 659303
rect 133081 659165 137580 659175
rect 5073 659093 14624 659103
rect 66170 659137 68582 659147
rect 5073 658727 14155 659093
rect 2509 658656 14155 658727
rect 79848 658972 82308 658982
rect 133210 658887 137580 659165
rect 139946 658887 140004 659558
rect 157083 659462 198006 659472
rect 133210 658850 140004 658887
rect 206714 659015 212383 659085
rect 206714 658768 209986 659015
rect 206585 658758 209986 658768
rect 206858 658630 209986 658758
rect 206585 658620 209986 658630
rect 79848 657975 82308 657985
rect 149997 658524 152333 658534
rect 66170 657860 68582 657870
rect 21160 657690 23631 657700
rect 23631 657665 23640 657675
rect 21160 657522 23640 657532
rect 124336 657669 126700 657679
rect 124336 657519 126700 657529
rect 206714 658377 209986 658620
rect 212293 658377 212383 659015
rect 206714 658305 212383 658377
rect 149997 657385 152333 657395
rect 34979 657242 35060 657252
rect 32682 657177 34979 657233
rect 34979 657153 35060 657163
rect 112670 657243 112802 657253
rect 112802 657177 115172 657233
rect 112670 657150 112802 657160
rect 197714 657125 199942 657135
rect 73065 657028 74069 657038
rect 34974 656786 35066 656796
rect 35452 656766 73065 656798
rect 35066 656710 73065 656766
rect 34974 656670 35066 656680
rect 35452 656678 73065 656710
rect 197714 656991 199942 657001
rect 186140 656702 186225 656712
rect 186225 656635 188420 656691
rect 186140 656613 186225 656623
rect 112636 656533 112797 656543
rect 74069 656363 112636 656488
rect 112636 656338 112797 656348
rect 152623 656403 186037 656431
rect 152623 656300 152633 656403
rect 73065 656212 74069 656222
rect 153791 656393 186037 656403
rect 186129 656414 186241 656424
rect 153791 656337 186129 656393
rect 153791 656300 186037 656337
rect 186129 656306 186241 656316
rect 152633 656124 153791 656134
rect 144160 637403 145498 637413
rect 125227 637291 144160 637369
rect 124857 637281 144160 637291
rect 125442 637057 144160 637281
rect 124857 637047 144160 637057
rect 125227 636972 144160 637047
rect 145498 636972 145544 637369
rect 144160 636927 145498 636937
rect 368681 635516 368816 635526
rect 368681 635411 368816 635421
rect 368680 633678 368815 633688
rect 368680 633573 368815 633583
rect 152624 510676 153820 510686
rect 1323 510540 152624 510561
rect 1323 510538 73012 510540
rect 1323 510236 1358 510538
rect 2171 510260 73012 510538
rect 74070 510260 152624 510540
rect 2171 510236 152624 510260
rect 1323 510212 152624 510236
rect 153820 510212 153853 510561
rect 152624 510195 153820 510205
rect 1326 467320 145524 467339
rect 1326 467316 144170 467320
rect 1326 467014 1361 467316
rect 2174 467014 144170 467316
rect 1326 467013 144170 467014
rect 145472 467013 145524 467320
rect 1326 466990 145524 467013
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 198295 687830 199269 688219
rect 207123 688222 210596 688623
rect 207123 687795 210595 688222
rect 210595 687795 210596 688222
rect 211169 688246 214642 688703
rect 227277 688273 230750 688664
rect 211169 687875 211176 688246
rect 211176 687875 214642 688246
rect 223060 687834 226864 688186
rect 227277 687846 230749 688273
rect 230749 687846 230750 688273
rect 227277 687836 230750 687846
rect 231330 688282 234803 688683
rect 231330 687855 234802 688282
rect 234802 687855 234803 688282
rect 235312 688292 238785 688693
rect 235312 687865 238784 688292
rect 238784 687865 238785 688292
rect 239333 688287 242806 688688
rect 239333 687860 242805 688287
rect 242805 687860 242806 688287
rect 243372 688285 246845 688686
rect 243372 687858 246844 688285
rect 246844 687858 246845 688285
rect 202780 685044 247142 685291
rect 202780 684711 247142 685044
rect 23042 660431 64025 660657
rect 23042 660101 64025 660431
rect 83765 660472 124085 660846
rect 83765 660179 112324 660472
rect 112324 660445 124085 660472
rect 112324 660332 120252 660445
rect 112324 660179 112657 660332
rect 112657 660179 119074 660332
rect 119074 660179 120252 660332
rect 120252 660179 124085 660445
rect 157083 659901 197708 660502
rect 2671 658727 5073 659760
rect 66170 657870 68582 659137
rect 79848 657985 82308 658972
rect 137580 658887 139946 659558
rect 157083 659472 197708 659901
rect 21160 657665 23631 657690
rect 21160 657532 23631 657665
rect 124336 657529 126700 657669
rect 149997 657395 152333 658524
rect 209986 658377 212293 659015
rect 73065 656222 74069 657028
rect 197714 657001 199942 657125
rect 152633 656134 153791 656403
rect 144160 636937 145498 637403
rect 368681 635421 368816 635516
rect 368680 633583 368815 633678
rect 1358 510236 2171 510538
rect 73012 510260 74070 510540
rect 152624 510205 153820 510676
rect 1361 467014 2174 467316
rect 144170 467013 145472 467320
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 703099 515394 704800
rect 520594 703099 525394 704800
rect 17496 693341 19996 702300
rect 69842 699968 72342 702300
rect 69842 697468 82326 699968
rect 17498 693242 19996 693341
rect 17498 690824 17558 693242
rect 19943 690824 19996 693242
rect 17498 690746 19996 690824
rect 66130 693229 68630 693269
rect 66130 690828 66188 693229
rect 68553 690828 68630 693229
rect -800 683796 1700 685242
rect -800 681296 5105 683796
rect 21882 681701 21892 683906
rect 22854 681701 22864 683906
rect -800 680242 1700 681296
rect 2605 659760 5105 681296
rect 2605 658727 2671 659760
rect 5073 658727 5105 659760
rect -800 643842 1660 648642
rect -800 633842 1660 638642
rect 2605 611726 5105 658727
rect 21889 657695 22824 681701
rect 23032 660101 23042 661269
rect 64017 660662 64027 661269
rect 64017 660657 64035 660662
rect 64025 660101 64035 660657
rect 23032 660096 64035 660101
rect 66130 659137 68630 690828
rect 66130 657870 66170 659137
rect 68582 657870 68630 659137
rect 79826 658972 82326 697468
rect 121407 699624 123907 702300
rect 121407 697124 152455 699624
rect 93805 695867 95820 695904
rect 93805 693909 93859 695867
rect 95764 693909 95820 695867
rect 93805 683893 95820 693909
rect 124995 692109 125005 692310
rect 93805 681853 93843 683893
rect 93833 681797 93843 681853
rect 95721 681853 95820 683893
rect 124989 690355 125005 692109
rect 125955 690355 125965 692310
rect 95721 681797 95731 681853
rect 83755 660179 83765 661487
rect 124071 660851 124081 661487
rect 124071 660846 124095 660851
rect 124085 660179 124095 660846
rect 83755 660174 124095 660179
rect 79826 657985 79848 658972
rect 82308 657985 82326 658972
rect 79826 657959 82326 657985
rect 21150 657690 23641 657695
rect 21150 657532 21160 657690
rect 23631 657532 23641 657690
rect 66130 657635 68630 657870
rect 124989 657674 125924 690355
rect 137480 659558 139980 659593
rect 137480 658887 137580 659558
rect 139946 658887 139980 659558
rect 124326 657669 126710 657674
rect 21150 657527 23641 657532
rect 124326 657529 124336 657669
rect 126700 657529 126710 657669
rect 124326 657524 126710 657529
rect 72999 657028 74122 657160
rect 72999 656222 73065 657028
rect 74069 656222 74122 657028
rect 14417 621627 14427 624619
rect 64644 621627 64654 624619
rect 2605 607134 2646 611726
rect 2636 607093 2646 607134
rect 5007 607134 5105 611726
rect 5007 607093 5017 607134
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect -800 511530 480 511642
rect 1348 510538 2181 510543
rect 1348 510460 1358 510538
rect -800 510348 1358 510460
rect 1292 510340 1358 510348
rect 1348 510236 1358 510340
rect 2171 510236 2181 510538
rect 1348 510231 2181 510236
rect 72999 510540 74122 656222
rect 83142 622007 83152 624630
rect 133410 622007 133420 624630
rect 137480 611839 139980 658887
rect 149955 658524 152455 697124
rect 166763 695391 169263 702300
rect 177015 695391 179515 702300
rect 218640 697309 221140 702300
rect 166762 692889 179515 695391
rect 211648 693981 211658 695778
rect 214091 695500 214101 695778
rect 214091 693981 214151 695500
rect 218640 694902 218717 697309
rect 221066 694902 221140 697309
rect 218640 694879 221140 694902
rect 223860 697338 226360 697368
rect 223860 694931 223921 697338
rect 226270 694931 226360 697338
rect 171983 684070 174483 692889
rect 207536 692355 210036 692388
rect 207536 690328 207591 692355
rect 209950 690328 210036 692355
rect 207536 688628 210036 690328
rect 211651 688708 214151 693981
rect 211159 688703 214652 688708
rect 207113 688623 210606 688628
rect 198292 688224 199274 688239
rect 198285 688219 199279 688224
rect 198285 687830 198295 688219
rect 199269 687830 199279 688219
rect 198285 687825 199279 687830
rect 171983 681570 192882 684070
rect 190382 667305 192882 681570
rect 190367 664796 190377 667305
rect 192874 664796 192884 667305
rect 157073 660502 197718 660507
rect 157073 659472 157083 660502
rect 197708 659472 197718 660502
rect 157073 659467 197718 659472
rect 149955 657395 149997 658524
rect 152333 657395 152455 658524
rect 149955 657301 152455 657395
rect 198292 657130 199274 687825
rect 207113 687795 207123 688623
rect 210596 687795 210606 688623
rect 211159 687875 211169 688703
rect 214642 687875 214652 688703
rect 223860 688191 226360 694931
rect 228892 697352 231392 702300
rect 242722 699634 242732 702134
rect 245232 702114 245242 702134
rect 245232 699634 315546 702114
rect 243372 699614 315546 699634
rect 228892 694945 228965 697352
rect 231314 694945 231392 697352
rect 228892 694833 231392 694945
rect 232116 696758 311894 699258
rect 232116 688688 234616 696758
rect 235915 693974 307678 696474
rect 235915 688698 238415 693974
rect 239738 691142 303725 693642
rect 235302 688693 238795 688698
rect 239738 688693 242238 691142
rect 231320 688683 234813 688688
rect 227267 688664 230760 688669
rect 211159 687870 214652 687875
rect 223050 688186 226874 688191
rect 223050 687834 223060 688186
rect 226864 687834 226874 688186
rect 223050 687829 226874 687834
rect 227267 687836 227277 688664
rect 230750 687836 230760 688664
rect 231320 687855 231330 688683
rect 234803 687855 234813 688683
rect 235302 687865 235312 688693
rect 238785 687865 238795 688693
rect 235302 687860 238795 687865
rect 239323 688688 242816 688693
rect 239323 687860 239333 688688
rect 242806 687860 242816 688688
rect 239323 687855 242816 687860
rect 243362 688686 299390 690785
rect 243362 687858 243372 688686
rect 246845 688285 299390 688686
rect 246845 687858 246855 688285
rect 231320 687850 234813 687855
rect 243362 687853 246855 687858
rect 227267 687831 230760 687836
rect 207113 687790 210606 687795
rect 202770 685291 247152 685296
rect 202770 684711 202780 685291
rect 247142 684711 247152 685291
rect 202770 684706 202805 684711
rect 202795 684082 202805 684706
rect 247109 684706 247152 684711
rect 247109 684082 247119 684706
rect 209899 659015 212399 659121
rect 209899 658377 209986 659015
rect 212293 658377 212399 659015
rect 197704 657125 199952 657130
rect 197704 657001 197714 657125
rect 199942 657001 199952 657125
rect 197704 656996 199952 657001
rect 152609 656403 153837 656431
rect 152609 656134 152633 656403
rect 153791 656134 153837 656403
rect 137480 607168 137755 611839
rect 139770 607168 139980 611839
rect 137480 607076 139980 607168
rect 144145 637403 145521 637418
rect 144145 636937 144160 637403
rect 145498 636937 145521 637403
rect 72999 510260 73012 510540
rect 74070 510260 74122 510540
rect 72999 510192 74122 510260
rect -800 509166 480 509278
rect -800 507984 490 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect 1351 467316 2184 467321
rect -800 467230 480 467238
rect 1351 467230 1361 467316
rect -800 467126 1361 467230
rect 304 467118 1361 467126
rect 1351 467014 1361 467118
rect 2174 467014 2184 467316
rect 1351 467009 2184 467014
rect 144145 467320 145521 636937
rect 152609 510676 153837 656134
rect 156490 620709 156500 624128
rect 206836 620709 206846 624128
rect 209899 611733 212399 658377
rect 296890 658340 299390 688285
rect 301225 661655 303725 691142
rect 305178 664670 307678 693974
rect 309394 668158 311894 696758
rect 313046 671728 315546 699614
rect 320335 695123 322835 702300
rect 330587 695123 333087 702300
rect 414564 696421 417064 702300
rect 466720 696421 469220 702300
rect 510501 696878 510511 703099
rect 525661 696878 525671 703099
rect 566594 702300 571594 704800
rect 567875 698736 570375 702300
rect 567865 696717 567875 698736
rect 570375 696717 570385 698736
rect 320334 692621 333087 695123
rect 414554 693921 414564 696421
rect 417064 693921 417074 696421
rect 466710 693921 466720 696421
rect 469220 693921 469230 696421
rect 313036 669228 313046 671728
rect 315546 669228 315556 671728
rect 309384 665658 309394 668158
rect 311894 665658 311904 668158
rect 305168 662170 305178 664670
rect 307678 662170 307688 664670
rect 301215 659155 301225 661655
rect 303725 659155 303735 661655
rect 296880 655840 296890 658340
rect 299390 655840 299400 658340
rect 325555 650863 328055 692621
rect 582300 681668 584800 682984
rect 576277 679168 576287 681668
rect 578306 679168 584800 681668
rect 582300 677984 584800 679168
rect 373465 669228 373475 671728
rect 374825 669228 374835 671728
rect 371778 665658 371788 668158
rect 373138 665658 373148 668158
rect 369963 662170 369973 664670
rect 371323 662170 371333 664670
rect 368199 661655 369549 661704
rect 368189 659155 368199 661655
rect 369549 659155 369559 661655
rect 366150 655840 366160 658340
rect 367510 655840 367520 658340
rect 325545 648363 325555 650863
rect 328055 648363 328065 650863
rect 325555 648358 328055 648363
rect 366160 642905 367510 655840
rect 368199 642905 369549 659155
rect 369973 642905 371323 662170
rect 371788 642905 373138 665658
rect 373475 642905 374825 669228
rect 367006 642208 367202 642905
rect 360862 642012 367202 642208
rect 347630 636697 347636 637147
rect 348086 636697 348966 637147
rect 360862 636883 361058 642012
rect 368630 641752 368826 642905
rect 368630 641556 370520 641752
rect 368671 635516 368826 635521
rect 368671 635421 368681 635516
rect 368816 635421 368826 635516
rect 368671 635418 368826 635421
rect 368652 635049 368848 635418
rect 370324 635049 370520 641556
rect 368652 634853 370520 635049
rect 370918 634243 371114 642905
rect 372372 642103 372568 642905
rect 371439 641907 372568 642103
rect 371439 637006 371635 641907
rect 374402 641653 374598 642905
rect 371879 641457 374598 641653
rect 368651 634047 371114 634243
rect 368651 633678 368847 634047
rect 368651 633588 368680 633678
rect 368670 633583 368680 633588
rect 368815 633588 368847 633678
rect 368815 633583 368825 633588
rect 368670 633578 368825 633583
rect 371879 632836 372075 641457
rect 582340 639784 584800 644584
rect 371440 632640 372075 632836
rect 371440 632181 371636 632640
rect 352226 630044 352236 630281
rect 352702 630044 352712 630281
rect 352226 613751 352712 630044
rect 356365 630025 356375 630262
rect 356841 630025 356851 630262
rect 356365 615037 356851 630025
rect 358816 630047 358826 630284
rect 359292 630047 359302 630284
rect 358816 616322 359302 630047
rect 582340 629784 584800 634584
rect 361089 628771 361575 628785
rect 360254 628619 360264 628648
rect 360218 628346 360264 628619
rect 360662 628619 360672 628648
rect 360662 628346 360704 628619
rect 360218 618008 360704 628346
rect 361089 628469 361132 628771
rect 361530 628469 361575 628771
rect 361089 619534 361575 628469
rect 362010 628738 362496 628770
rect 362010 628436 362048 628738
rect 362446 628436 362496 628738
rect 362010 620980 362496 628436
rect 362010 620494 383337 620980
rect 382851 619658 383337 620494
rect 361089 619048 379241 619534
rect 360218 617522 374744 618008
rect 378755 617971 379241 619048
rect 374258 616445 374744 617522
rect 358816 615836 369845 616322
rect 356365 614551 365990 615037
rect 369359 614999 369845 615836
rect 352226 613265 360609 613751
rect 360123 612028 360609 613265
rect 365504 613072 365990 614551
rect 209899 607161 210137 611733
rect 212245 607161 212399 611733
rect 209899 606979 212399 607161
rect 152609 510205 152624 510676
rect 153820 510205 153837 510676
rect 152609 510169 153837 510205
rect 144145 467013 144170 467320
rect 145472 467013 145521 467320
rect 144145 466948 145521 467013
rect -800 465944 480 466056
rect -800 464872 1188 464874
rect -800 464762 1508 464872
rect 253 464760 1508 464762
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 359161 315293 361661 612028
rect 363819 361386 366319 613072
rect 368397 407710 370897 614999
rect 373136 452031 375636 616445
rect 377553 496436 380053 617971
rect 381890 581162 384390 619658
rect 583554 589472 584800 589584
rect 583554 588290 584800 588402
rect 583554 587108 584800 587220
rect 583554 585926 584800 586038
rect 570571 584856 580767 585210
rect 570571 584744 584800 584856
rect 570571 582710 580767 584744
rect 583554 583562 584800 583674
rect 570571 581162 573071 582710
rect 381890 578662 573071 581162
rect 578758 540186 578768 555678
rect 583178 555362 583188 555678
rect 583178 550562 584800 555362
rect 583178 545362 583188 550562
rect 583178 540562 584800 545362
rect 583178 540186 583188 540562
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 377553 495434 581308 496436
rect 377553 495322 584800 495434
rect 377553 493936 581308 495322
rect 583520 494140 584800 494252
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 373136 451012 581762 452031
rect 373136 450900 584800 451012
rect 373136 449531 581762 450900
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 368397 406590 581354 407710
rect 583520 407660 584800 407772
rect 368397 406478 584800 406590
rect 368397 405210 581354 406478
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 363819 360168 580825 361386
rect 583520 361238 584800 361350
rect 363819 360056 584800 360168
rect 363819 358886 580825 360056
rect 583520 358874 584800 358986
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 359161 314946 581320 315293
rect 359161 314834 584800 314946
rect 359161 312793 581320 314834
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 578927 240347 581622 240589
rect 578409 225380 578419 240347
rect 583286 240030 583296 240347
rect 583286 235230 584800 240030
rect 583286 230030 583296 235230
rect 583286 225380 584800 230030
rect 578927 225230 584800 225380
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 151577 584800 151630
rect 578897 136610 578907 151577
rect 583774 146830 584800 151577
rect 583774 141630 583784 146830
rect 583774 136830 584800 141630
rect 583774 136610 583784 136830
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 17558 690824 19943 693242
rect 66188 690828 68553 693229
rect 21892 681701 22854 683906
rect 23042 660657 64017 661269
rect 23042 660101 64017 660657
rect 93859 693909 95764 695867
rect 93843 681797 95721 683893
rect 125005 690355 125955 692310
rect 83765 660846 124071 661487
rect 83765 660179 124071 660846
rect 14427 621627 64644 624619
rect 2646 607093 5007 611726
rect 83152 622007 133410 624630
rect 211658 693981 214091 695778
rect 218717 694902 221066 697309
rect 223921 694931 226270 697338
rect 207591 690328 209950 692355
rect 190377 664796 192874 667305
rect 157083 659472 197708 660502
rect 242732 699634 245232 702134
rect 228965 694945 231314 697352
rect 227277 688115 230750 688664
rect 202780 684711 247142 685291
rect 202805 684082 247109 684711
rect 137755 607168 139770 611839
rect 156500 620709 206836 624128
rect 510511 696878 525661 703099
rect 567875 696717 570375 698736
rect 414564 693921 417064 696421
rect 466720 693921 469220 696421
rect 313046 669228 315546 671728
rect 309394 665658 311894 668158
rect 305178 662170 307678 664670
rect 301225 659155 303725 661655
rect 296890 655840 299390 658340
rect 576287 679168 578306 681668
rect 373475 669228 374825 671728
rect 371788 665658 373138 668158
rect 369973 662170 371323 664670
rect 368199 659155 369549 661655
rect 366160 655840 367510 658340
rect 325555 648363 328055 650863
rect 347636 636697 348086 637147
rect 352236 630044 352702 630281
rect 356375 630025 356841 630262
rect 358826 630047 359292 630284
rect 360264 628346 360662 628648
rect 361132 628469 361530 628771
rect 362048 628436 362446 628738
rect 210137 607161 212245 611733
rect 578768 540186 583178 555678
rect 578419 225380 583286 240347
rect 578907 136610 583774 151577
<< metal4 >>
rect 510510 703099 525662 703100
rect 242731 702134 245233 702135
rect 242731 699634 242732 702134
rect 245232 699634 245233 702134
rect 242731 699633 245233 699634
rect 218687 697352 231368 697368
rect 218687 697338 228965 697352
rect 218687 697309 223921 697338
rect 93805 695867 214125 695904
rect 93805 693909 93859 695867
rect 95764 695778 214125 695867
rect 95764 693981 211658 695778
rect 214091 693981 214125 695778
rect 218687 694902 218717 697309
rect 221066 694931 223921 697309
rect 226270 694945 228965 697338
rect 231314 694945 231368 697352
rect 510510 696878 510511 703099
rect 525661 696878 525662 703099
rect 510510 696877 525662 696878
rect 567874 698736 570376 698737
rect 567874 696717 567875 698736
rect 570375 696717 570376 698736
rect 567874 696716 570376 696717
rect 226270 694931 231368 694945
rect 221066 694902 231368 694931
rect 218687 694868 231368 694902
rect 414563 696421 417065 696422
rect 95764 693909 214125 693981
rect 414563 693921 414564 696421
rect 417064 693921 417065 696421
rect 414563 693920 417065 693921
rect 466719 696421 469221 696422
rect 466719 693921 466720 696421
rect 469220 693921 469221 696421
rect 466719 693920 469221 693921
rect 93805 693889 214125 693909
rect 17498 693242 68630 693269
rect 17498 690824 17558 693242
rect 19943 693229 68630 693242
rect 19943 690828 66188 693229
rect 68553 690828 68630 693229
rect 207590 692355 209951 692356
rect 207590 692349 207591 692355
rect 19943 690824 68630 690828
rect 17498 690769 68630 690824
rect 124977 692310 207591 692349
rect 124977 690355 125005 692310
rect 125955 690355 207591 692310
rect 124977 690334 207591 690355
rect 207590 690328 207591 690334
rect 209950 690328 209951 692355
rect 207590 690327 209951 690328
rect 567875 690311 570375 696716
rect 227276 688664 230751 688665
rect 227276 688115 227277 688664
rect 230750 688115 230751 688664
rect 227276 688114 230751 688115
rect 536686 687811 570375 690311
rect 202779 685291 247143 685292
rect 202779 685235 202780 685291
rect 247142 684711 247143 685291
rect 247109 684710 247143 684711
rect 21910 683907 95867 683939
rect 21891 683906 95867 683907
rect 21891 681701 21892 683906
rect 22854 683893 95867 683906
rect 22854 681797 93843 683893
rect 95721 681797 95867 683893
rect 247109 684081 247110 684710
rect 22854 681710 95867 681797
rect 22854 681701 22855 681710
rect 21891 681700 22855 681701
rect 31160 677876 260437 677902
rect 31160 677857 142936 677876
rect 31160 677668 72143 677857
rect 46493 673154 72143 677668
rect 31160 673096 72143 673154
rect 75277 677786 142936 677857
rect 75277 673232 101968 677786
rect 117567 673232 142936 677786
rect 75277 673096 142936 673232
rect 31160 673047 142936 673096
rect 145430 677841 260437 677876
rect 145430 677818 216578 677841
rect 145430 673110 171320 677818
rect 184865 673110 216578 677818
rect 145430 673047 216578 673110
rect 31160 673035 216578 673047
rect 232215 673035 260437 677841
rect 274962 677887 467817 677902
rect 274962 673047 452327 677887
rect 467023 673047 467817 677887
rect 274962 673035 467817 673047
rect 313045 671728 315547 671729
rect 373474 671728 374826 671729
rect 313045 669228 313046 671728
rect 315546 669228 373475 671728
rect 374825 669228 374835 671728
rect 313045 669227 315547 669228
rect 373474 669227 374826 669228
rect 309393 668158 311895 668159
rect 371787 668158 373139 668159
rect 190376 667305 192875 667306
rect 190376 664796 190377 667305
rect 192874 667299 192875 667305
rect 192874 664799 235517 667299
rect 309393 665658 309394 668158
rect 311894 665658 371788 668158
rect 373138 665658 373148 668158
rect 309393 665657 311895 665658
rect 371787 665657 373139 665658
rect 192874 664796 192875 664799
rect 190376 664795 192875 664796
rect 23041 660101 23042 661270
rect 64017 660101 64018 661270
rect 83764 660179 83765 661488
rect 83764 660178 124072 660179
rect 23041 660100 64018 660101
rect 157082 659472 157083 660503
rect 197702 660502 197709 660503
rect 197708 659472 197709 660502
rect 157082 659471 197709 659472
rect 233017 635570 235517 664799
rect 305177 664670 307679 664671
rect 369972 664670 371324 664671
rect 305177 662170 305178 664670
rect 307678 662170 369973 664670
rect 371323 662170 371333 664670
rect 305177 662169 307679 662170
rect 369972 662169 371324 662170
rect 301224 661655 303726 661656
rect 368198 661655 369550 661656
rect 301224 659155 301225 661655
rect 303725 659155 368199 661655
rect 369549 659155 369559 661655
rect 301224 659154 303726 659155
rect 368198 659154 369550 659155
rect 296889 658340 299391 658341
rect 366159 658340 367511 658341
rect 296889 655840 296890 658340
rect 299390 655840 366160 658340
rect 367510 655840 367520 658340
rect 296889 655839 299391 655840
rect 366159 655839 367511 655840
rect 325554 650863 328056 650864
rect 251036 648363 325555 650863
rect 328055 648363 328065 650863
rect 251036 643769 253536 648363
rect 325554 648362 328056 648363
rect 251036 641269 338266 643769
rect 356990 643636 357847 643763
rect 357720 642897 357847 643636
rect 358200 643636 359056 643763
rect 358200 642897 358327 643636
rect 335766 640142 338266 641269
rect 335766 639692 348716 640142
rect 536686 639819 539186 687811
rect 576286 681668 578307 681669
rect 383342 637319 539186 639819
rect 544840 679168 576287 681668
rect 578306 679168 578307 681668
rect 347635 637147 348087 637148
rect 335766 636697 347636 637147
rect 348086 636697 348087 637147
rect 335766 635570 338266 636697
rect 347635 636696 348087 636697
rect 383342 635788 383892 637319
rect 376970 635579 383892 635788
rect 233017 633070 338266 635570
rect 376994 633304 383892 633513
rect 352335 630282 352605 632949
rect 352235 630281 352703 630282
rect 352235 630044 352236 630281
rect 352702 630044 352703 630281
rect 356477 630263 356747 632977
rect 358930 630285 359200 632879
rect 383342 631773 383892 633304
rect 544840 631773 547340 679168
rect 576286 679167 578307 679168
rect 358825 630284 359293 630285
rect 352235 630043 352703 630044
rect 356374 630262 356842 630263
rect 356374 630025 356375 630262
rect 356841 630025 356842 630262
rect 358825 630047 358826 630284
rect 359292 630047 359293 630284
rect 358825 630046 359293 630047
rect 356374 630024 356842 630025
rect 383342 629273 547340 631773
rect 361131 628771 361531 628772
rect 360263 628648 360663 628649
rect 360263 628346 360264 628648
rect 360662 628346 360663 628648
rect 361131 628469 361132 628771
rect 361530 628469 361531 628771
rect 361131 628468 361531 628469
rect 362047 628738 362447 628739
rect 362047 628436 362048 628738
rect 362446 628436 362447 628738
rect 362047 628435 362447 628436
rect 360263 628345 360663 628346
rect 14426 624619 64645 624620
rect 14426 624437 14427 624619
rect 64644 621627 64645 624619
rect 64282 621626 64645 621627
rect 156499 624128 206837 624129
rect 156499 624087 156500 624128
rect 206836 620708 206837 624128
rect 275302 624644 345528 625028
rect 275302 617580 311280 624644
rect 345358 623908 345528 624644
rect 345358 621915 380146 623908
rect 345358 617580 345528 621915
rect 275302 617272 345528 617580
rect 2575 611839 212044 611907
rect 2575 611726 137755 611839
rect 2575 607093 2646 611726
rect 5007 607168 137755 611726
rect 139770 611734 212044 611839
rect 139770 611733 212246 611734
rect 139770 607168 210137 611733
rect 5007 607161 210137 607168
rect 212245 607161 212246 611733
rect 5007 607160 212246 607161
rect 5007 607093 212044 607160
rect 2575 607040 212044 607093
rect 30038 599282 561785 599316
rect 30038 583701 30180 599282
rect 46130 599210 561785 599282
rect 46130 599176 147711 599210
rect 151098 599184 561785 599210
rect 151098 599176 381126 599184
rect 46130 599172 124862 599176
rect 46130 599145 51929 599172
rect 67434 599127 124862 599172
rect 30038 583663 41447 583701
rect 67434 583668 77083 599127
rect 67237 583663 77083 583668
rect 30038 583498 77083 583663
rect 79747 598859 124862 599127
rect 79747 583498 100668 598859
rect 30038 583445 100668 583498
rect 116512 583547 124862 598859
rect 154759 599126 381126 599176
rect 154759 599018 289653 599126
rect 154759 598949 195851 599018
rect 154759 583674 172469 598949
rect 187791 583729 195851 598949
rect 227970 583729 289653 599018
rect 187791 583674 289653 583729
rect 154759 583547 289653 583674
rect 116512 583507 147711 583547
rect 151098 583507 289653 583547
rect 116512 583497 289653 583507
rect 319550 598747 381126 599126
rect 319550 583865 338602 598747
rect 353942 583865 381126 598747
rect 319550 583555 381126 583865
rect 411023 599165 561785 599184
rect 411023 583555 487932 599165
rect 319550 583536 487932 583555
rect 525630 598800 561785 599165
rect 525630 584066 546176 598800
rect 561217 584066 561785 598800
rect 525630 583536 561785 584066
rect 319550 583497 561785 583536
rect 116512 583445 561785 583497
rect 20619 555772 583382 555900
rect 32921 555678 583382 555772
rect 32921 555640 578768 555678
rect 32921 555464 259862 555640
rect 32921 555414 199695 555464
rect 32921 540298 40996 555414
rect 70830 555351 199695 555414
rect 70830 540407 128975 555351
rect 159252 540409 199695 555351
rect 229967 540435 259862 555464
rect 275226 555601 578768 555640
rect 275226 555588 452164 555601
rect 275226 555313 385148 555588
rect 275226 540435 293791 555313
rect 229967 540409 293791 540435
rect 159252 540407 293791 540409
rect 70830 540369 293791 540407
rect 324068 540644 385148 555313
rect 415425 540644 452164 555588
rect 324068 540369 452164 540644
rect 70830 540298 452164 540369
rect 32921 540202 452164 540298
rect 20619 540149 452164 540202
rect 467493 555349 578768 555601
rect 467493 540466 491313 555349
rect 521955 540466 578768 555349
rect 467493 540186 578768 540466
rect 583178 540186 583382 555678
rect 467493 540149 583382 540186
rect 20619 540029 583382 540149
rect 102586 432559 557291 432965
rect 102586 432558 338894 432559
rect 116402 417742 338894 432558
rect 354227 432093 557291 432559
rect 354227 417742 545705 432093
rect 116402 417422 545705 417742
rect 102586 417276 545705 417422
rect 102586 417094 557291 417276
rect 21612 378918 466454 379014
rect 21612 378759 452093 378918
rect 21612 378616 259965 378759
rect 33021 363349 259965 378616
rect 21612 363295 259965 363349
rect 275183 363464 452093 378759
rect 275183 363295 466454 363464
rect 21612 363143 466454 363295
rect 22911 240605 583795 240685
rect 32695 240427 583795 240605
rect 32695 225260 259755 240427
rect 275011 240355 583795 240427
rect 275011 225376 452031 240355
rect 467535 240347 583795 240355
rect 467535 225380 578419 240347
rect 583286 225380 583795 240347
rect 467535 225376 583795 225380
rect 275011 225260 583795 225376
rect 32695 225102 583795 225260
rect 22911 225078 583795 225102
rect 563330 225074 578151 225078
rect 100326 151702 583784 151892
rect 100326 151653 545482 151702
rect 100326 151638 338641 151653
rect 100326 136586 100582 151638
rect 116556 136586 338641 151638
rect 100326 136461 338641 136586
rect 354383 136619 545482 151653
rect 561448 151577 583784 151702
rect 561448 136619 578907 151577
rect 354383 136610 578907 136619
rect 583774 136610 583784 151577
rect 354383 136461 583784 136610
rect 100326 136443 583784 136461
<< via4 >>
rect 242732 699634 245232 702134
rect 510511 696878 525661 703099
rect 414564 693921 417064 696421
rect 466720 693921 469220 696421
rect 227277 688115 230750 688664
rect 202733 684711 202780 685235
rect 202780 684711 247109 685235
rect 202733 684082 202805 684711
rect 202805 684082 247109 684711
rect 202733 683217 247109 684082
rect 31049 673154 46493 677668
rect 72143 673096 75277 677857
rect 101968 673232 117567 677786
rect 142936 673047 145430 677876
rect 171320 673110 184865 677818
rect 216578 672994 232215 677841
rect 260437 671893 274962 678175
rect 452327 673047 467023 677887
rect 23042 661269 64017 661882
rect 23042 660101 64017 661269
rect 83765 661487 124085 662834
rect 83765 660179 124071 661487
rect 124071 660179 124085 661487
rect 157083 660502 197702 661420
rect 157083 659472 197702 660502
rect 356670 643622 356990 643930
rect 359056 643622 359376 643930
rect 360315 637262 360607 637553
rect 361033 637228 361327 637566
rect 362102 637245 362396 637583
rect 360264 628346 360662 628648
rect 361132 628469 361530 628771
rect 362048 628436 362446 628738
rect 83049 624683 133410 624733
rect 82973 624630 133488 624683
rect 14337 621627 14427 624437
rect 14427 621627 64282 624437
rect 14337 618001 64282 621627
rect 82973 622007 83152 624630
rect 83152 622007 133410 624630
rect 133410 622007 133488 624630
rect 82973 617893 133488 622007
rect 156376 620709 156500 624087
rect 156500 620709 206836 624087
rect 156376 619144 206836 620709
rect 259670 617074 275302 625270
rect 311280 617580 345358 624644
rect 380146 621915 380589 623908
rect 30180 599145 46130 599282
rect 147711 599176 151098 599210
rect 51929 599145 67434 599172
rect 30180 583701 67434 599145
rect 41447 583668 67434 583701
rect 41447 583663 67237 583668
rect 77083 583498 79747 599127
rect 100668 583221 116512 598859
rect 124862 583547 154759 599176
rect 172469 583674 187791 598949
rect 195851 583729 227970 599018
rect 147711 583507 151098 583547
rect 289653 583497 319550 599126
rect 338602 583865 353942 598747
rect 381126 583555 411023 599184
rect 487932 583536 525630 599165
rect 546176 584066 561217 598800
rect 17921 540202 32921 555772
rect 40996 540298 70830 555414
rect 128975 540407 159252 555351
rect 199695 540409 229967 555464
rect 259862 540435 275226 555640
rect 293791 540369 324068 555313
rect 385148 540644 415425 555588
rect 452164 540149 467493 555601
rect 491313 540466 521955 555349
rect 101051 417422 116402 432558
rect 338894 417742 354227 432559
rect 545705 417276 561038 432093
rect 17721 363349 33021 378616
rect 259965 363295 275183 378759
rect 452093 363464 467213 378918
rect 17911 225102 32695 240605
rect 259755 225260 275011 240427
rect 452031 225376 467535 240355
rect 100582 136586 116556 151638
rect 338641 136461 354383 151653
rect 545482 136619 561448 151702
<< metal5 >>
rect 510306 703099 525839 703217
rect 242708 702134 245256 702158
rect 242708 699634 242732 702134
rect 245232 699634 245256 702134
rect 242708 699610 245256 699634
rect 242732 693377 245232 699610
rect 510306 696878 510511 703099
rect 525661 696878 525839 703099
rect 414540 696421 417088 696445
rect 466696 696421 469244 696445
rect 414540 693921 414564 696421
rect 417064 693921 436162 696421
rect 414540 693897 417088 693921
rect 227790 690877 245232 693377
rect 227790 688688 230290 690877
rect 433662 690218 436162 693921
rect 227253 688664 230774 688688
rect 227253 688115 227277 688664
rect 230750 688115 230774 688664
rect 227253 688091 230774 688115
rect 352750 687718 436162 690218
rect 441224 693921 466720 696421
rect 469220 693921 469244 696421
rect 202709 685235 247133 685259
rect 202709 683217 202733 685235
rect 247109 683217 247133 685235
rect 202709 683193 247133 683217
rect 30960 677668 46833 678350
rect 30960 673154 31049 677668
rect 46493 673154 46833 677668
rect 30960 661906 46833 673154
rect 72119 677857 75301 677881
rect 72119 673096 72143 677857
rect 75277 677536 75301 677857
rect 142912 677876 145454 677900
rect 101944 677786 117591 677810
rect 75277 673096 75313 677536
rect 101944 677524 101968 677786
rect 72119 673072 75313 673096
rect 23018 661882 64041 661906
rect 23018 660101 23042 661882
rect 64017 660101 64041 661882
rect 23018 660077 64041 660101
rect 14313 624437 64306 624461
rect 14313 618001 14337 624437
rect 64282 618001 64306 624437
rect 14313 617977 64306 618001
rect 30017 599282 46173 617977
rect 72165 615148 75313 673072
rect 101864 673232 101968 677524
rect 117567 677524 117591 677786
rect 142912 677705 142936 677876
rect 117567 673232 117672 677524
rect 77216 613098 79845 671573
rect 101864 662858 117672 673232
rect 142885 673047 142936 677705
rect 145430 677705 145454 677876
rect 216581 677865 232247 683193
rect 171296 677818 184889 677842
rect 145430 673047 145500 677705
rect 171296 677636 171320 677818
rect 83741 662834 124109 662858
rect 83741 660179 83765 662834
rect 124085 660179 124109 662834
rect 83741 660155 124109 660179
rect 83025 624733 133434 624757
rect 83025 624707 83049 624733
rect 82949 624683 83049 624707
rect 133410 624707 133434 624733
rect 133410 624683 133512 624707
rect 82949 617893 82973 624683
rect 133488 617893 133512 624683
rect 82949 617869 133512 617893
rect 30017 586019 30180 599282
rect 46130 599169 46173 599282
rect 51497 599196 53807 599338
rect 58426 599196 60736 599292
rect 65356 599196 67666 599323
rect 51497 599172 67666 599196
rect 51497 599169 51929 599172
rect 46130 599145 51929 599169
rect 30156 583701 30180 586019
rect 30156 583677 41447 583701
rect 36223 560658 38615 583677
rect 41423 583663 41447 583677
rect 67434 583668 67666 599172
rect 67237 583663 67666 583668
rect 41423 583639 67666 583663
rect 44501 581203 46811 583639
rect 51497 581259 53807 583639
rect 45425 580076 45745 581203
rect 52369 580076 52689 581259
rect 58426 581098 60736 583639
rect 65356 581205 67666 583639
rect 77058 599127 79845 613098
rect 77058 583524 77083 599127
rect 77059 583498 77083 583524
rect 79747 583612 79845 599127
rect 100463 598859 116619 617869
rect 142885 615246 145500 673047
rect 171295 673110 171320 677636
rect 184865 673110 184889 677818
rect 171295 673086 184889 673110
rect 216554 677841 232247 677865
rect 79747 583498 79771 583612
rect 77059 583474 79771 583498
rect 100463 583221 100668 598859
rect 116512 583221 116619 598859
rect 59313 580076 59633 581098
rect 66257 580076 66577 581205
rect 17569 555772 33235 556317
rect 17569 540202 17921 555772
rect 32921 540202 33235 555772
rect 17569 378616 33235 540202
rect 40864 555438 43451 578397
rect 48022 555438 50609 578656
rect 54834 555438 57421 578570
rect 61819 555438 64406 578052
rect 68545 555438 71132 578483
rect 40864 555414 71132 555438
rect 40864 540298 40996 555414
rect 70830 540298 71132 555414
rect 40864 540274 71132 540298
rect 40864 540137 43451 540274
rect 48022 540113 50609 540274
rect 54834 540113 57421 540274
rect 61819 540137 64406 540274
rect 68545 540212 71132 540274
rect 17569 363349 17721 378616
rect 33021 363349 33235 378616
rect 17569 240605 33235 363349
rect 17569 225102 17911 240605
rect 32695 225102 33235 240605
rect 17569 224794 33235 225102
rect 100463 432558 116619 583221
rect 124759 599200 126962 599322
rect 147647 599210 151189 672301
rect 171295 661444 184887 673086
rect 216554 672994 216578 677841
rect 232215 673051 232247 677841
rect 259666 678175 275332 678276
rect 232215 672994 232239 673051
rect 216554 672970 232239 672994
rect 157059 661420 197726 661444
rect 157059 659472 157083 661420
rect 197702 659472 197726 661420
rect 157059 659448 197726 659472
rect 156352 624096 206860 624111
rect 156352 624087 207124 624096
rect 156352 619144 156376 624087
rect 206836 619144 207124 624087
rect 156352 619120 207124 619144
rect 147647 599200 147711 599210
rect 124759 599176 147711 599200
rect 151098 599200 151189 599210
rect 154493 599200 154813 599217
rect 151098 599176 154813 599200
rect 124759 583547 124862 599176
rect 154759 583547 154813 599176
rect 172171 598949 188327 619120
rect 218723 615607 222084 672970
rect 259666 671893 260437 678175
rect 274962 671893 275332 678175
rect 223844 599042 227386 658283
rect 259666 625294 275332 671893
rect 352750 647598 355250 687718
rect 441224 684427 443724 693921
rect 466696 693897 469244 693921
rect 360796 681927 443724 684427
rect 360796 647598 363296 681927
rect 352750 647048 356990 647598
rect 356670 643954 356990 647048
rect 359056 647048 363296 647598
rect 451976 677887 467642 678029
rect 451976 673047 452327 677887
rect 467023 673047 467642 677887
rect 359056 643954 359376 647048
rect 356646 643930 357014 643954
rect 356646 643622 356670 643930
rect 356990 643622 357014 643930
rect 356646 643598 357014 643622
rect 359032 643930 359400 643954
rect 359032 643622 359056 643930
rect 359376 643622 359400 643930
rect 359032 643598 359400 643622
rect 360291 637553 360631 637577
rect 360291 637262 360315 637553
rect 360607 637427 360631 637553
rect 361009 637566 361351 637590
rect 360607 637262 360633 637427
rect 259646 625270 275332 625294
rect 259646 617074 259670 625270
rect 275302 617074 275332 625270
rect 344840 624668 345283 631382
rect 346785 627046 347228 631405
rect 360291 628672 360633 637262
rect 361009 637228 361033 637566
rect 361327 637228 361351 637566
rect 361009 636893 361351 637228
rect 362078 637583 362420 637607
rect 362078 637245 362102 637583
rect 362396 637245 362420 637583
rect 361009 628795 361344 636893
rect 361009 628771 361554 628795
rect 360240 628648 360686 628672
rect 360240 628346 360264 628648
rect 360662 628346 360686 628648
rect 361009 628473 361132 628771
rect 361108 628469 361132 628473
rect 361530 628469 361554 628771
rect 362078 628762 362420 637245
rect 361108 628445 361554 628469
rect 362024 628738 362470 628762
rect 362024 628436 362048 628738
rect 362446 628436 362470 628738
rect 362024 628412 362470 628436
rect 360240 628322 360686 628346
rect 378201 627046 378644 630294
rect 346785 625053 378644 627046
rect 311256 624644 345382 624668
rect 311256 617580 311280 624644
rect 345358 617580 345382 624644
rect 311256 617556 345382 617580
rect 259646 617050 275332 617074
rect 195827 599018 227994 599042
rect 195827 598960 195851 599018
rect 172171 583913 172469 598949
rect 172445 583674 172469 583913
rect 187791 583913 188327 598949
rect 187791 583674 187815 583913
rect 172445 583650 187815 583674
rect 195244 583729 195851 598960
rect 227970 583729 227994 599018
rect 195244 583705 227994 583729
rect 124759 583523 147711 583547
rect 124759 560338 126962 583523
rect 133661 579201 133981 583523
rect 140605 579201 140925 583523
rect 147549 583507 147711 583523
rect 151098 583523 154813 583547
rect 151098 583507 151122 583523
rect 147549 583483 151122 583507
rect 147549 578864 147869 583483
rect 154493 579201 154813 583523
rect 195244 579563 197447 583705
rect 195244 579361 197522 579563
rect 128823 555375 131710 577101
rect 135608 555375 138495 576885
rect 143114 555375 146001 576957
rect 149754 555375 152641 577029
rect 156683 555375 159570 576740
rect 195244 573243 197447 579361
rect 197480 573243 197522 579361
rect 204146 579361 204466 583705
rect 197842 579262 203810 579286
rect 197842 573342 197866 579262
rect 199308 573342 202195 577261
rect 203786 573342 203810 579262
rect 197842 573318 203810 573342
rect 195244 572839 197522 573243
rect 195244 566721 197447 572839
rect 197480 566721 197522 572839
rect 199308 572764 202195 573318
rect 204146 573243 204188 579361
rect 204424 573243 204466 579361
rect 211090 579361 211410 583705
rect 204786 579262 210754 579286
rect 204786 573342 204810 579262
rect 206093 573342 208980 577045
rect 210730 573342 210754 579262
rect 204786 573318 210754 573342
rect 204146 572839 204466 573243
rect 197842 572740 203810 572764
rect 197842 566820 197866 572740
rect 199308 566820 202195 572740
rect 203786 566820 203810 572740
rect 197842 566796 203810 566820
rect 195244 566317 197522 566721
rect 195244 560199 197447 566317
rect 197480 560199 197522 566317
rect 199308 566242 202195 566796
rect 204146 566721 204188 572839
rect 204424 566721 204466 572839
rect 206093 572764 208980 573318
rect 211090 573243 211132 579361
rect 211368 573243 211410 579361
rect 211730 579262 216581 579286
rect 211730 573342 211754 579262
rect 218034 579243 218354 583705
rect 224978 579243 225298 583705
rect 213599 573342 216486 577117
rect 211730 573318 216581 573342
rect 211090 572839 211410 573243
rect 204786 572740 210754 572764
rect 204786 566820 204810 572740
rect 206093 566820 208980 572740
rect 210730 566820 210754 572740
rect 204786 566796 210754 566820
rect 204146 566317 204466 566721
rect 197842 566218 203810 566242
rect 197842 560298 197866 566218
rect 199308 560298 202195 566218
rect 203786 560298 203810 566218
rect 197842 560274 203810 560298
rect 195244 560051 197522 560199
rect 197202 559997 197522 560051
rect 128823 555351 159570 555375
rect 128823 540407 128975 555351
rect 159252 540407 159570 555351
rect 199308 555488 202195 560274
rect 204146 560199 204188 566317
rect 204424 560199 204466 566317
rect 206093 566242 208980 566796
rect 211090 566721 211132 572839
rect 211368 566721 211410 572839
rect 213599 572764 216486 573318
rect 211730 572740 216581 572764
rect 211730 566820 211754 572740
rect 213599 566820 216486 572740
rect 211730 566796 216581 566820
rect 211090 566317 211410 566721
rect 204786 566218 210754 566242
rect 204786 560298 204810 566218
rect 206093 560298 208980 566218
rect 210730 560298 210754 566218
rect 204786 560274 210754 560298
rect 204146 559997 204466 560199
rect 206093 555488 208980 560274
rect 211090 560199 211132 566317
rect 211368 560199 211410 566317
rect 213599 566242 216486 566796
rect 211730 566218 216581 566242
rect 211730 560298 211754 566218
rect 213599 560298 216486 566218
rect 211730 560274 216581 560298
rect 211090 559997 211410 560199
rect 213599 555488 216486 560274
rect 220132 555488 223019 578371
rect 227397 555488 230284 578371
rect 199308 555464 230284 555488
rect 199308 540415 199695 555464
rect 128823 540383 159570 540407
rect 199671 540409 199695 540415
rect 229967 540415 230284 555464
rect 259666 555640 275332 617050
rect 312320 604344 315940 617556
rect 319399 604291 323019 617556
rect 326025 604364 329645 617556
rect 333307 604619 336927 617556
rect 340152 604546 343772 617556
rect 346785 615384 354541 625053
rect 380146 623932 380589 631171
rect 380122 623908 380613 623932
rect 380122 621915 380146 623908
rect 380589 621915 380613 623908
rect 380122 621891 380613 621915
rect 345371 602316 354541 615384
rect 317349 600961 317669 602316
rect 324293 600961 324613 602316
rect 331237 600961 331557 602316
rect 338181 600961 338501 602316
rect 345125 600961 354541 602316
rect 317349 600926 354541 600961
rect 289452 599150 291655 599152
rect 317078 599150 354541 600926
rect 289452 599126 354541 599150
rect 289452 583497 289653 599126
rect 319550 598747 354541 599126
rect 319550 598383 338602 598747
rect 319550 583497 319574 598383
rect 338578 597776 338602 598383
rect 289452 583473 319574 583497
rect 338385 583865 338602 597776
rect 353942 583865 354541 598747
rect 381102 599184 411047 599208
rect 381102 598681 381126 599184
rect 289452 579107 291655 583473
rect 289452 578905 291730 579107
rect 289452 572787 291655 578905
rect 291688 572787 291730 578905
rect 298354 578905 298674 583473
rect 292050 578806 298018 578830
rect 292050 572886 292074 578806
rect 293516 572886 296403 576805
rect 297994 572886 298018 578806
rect 292050 572862 298018 572886
rect 289452 572383 291730 572787
rect 289452 566265 291655 572383
rect 291688 566265 291730 572383
rect 293516 572308 296403 572862
rect 298354 572787 298396 578905
rect 298632 572787 298674 578905
rect 305298 578905 305618 583473
rect 298994 578806 304962 578830
rect 298994 572886 299018 578806
rect 300301 572886 303188 576589
rect 304938 572886 304962 578806
rect 298994 572862 304962 572886
rect 298354 572383 298674 572787
rect 292050 572284 298018 572308
rect 292050 566364 292074 572284
rect 293516 566364 296403 572284
rect 297994 566364 298018 572284
rect 292050 566340 298018 566364
rect 289452 565861 291730 566265
rect 289452 560042 291655 565861
rect 291410 559743 291452 560042
rect 291688 559743 291730 565861
rect 293516 565786 296403 566340
rect 298354 566265 298396 572383
rect 298632 566265 298674 572383
rect 300301 572308 303188 572862
rect 305298 572787 305340 578905
rect 305576 572787 305618 578905
rect 312242 578905 312562 583473
rect 305938 578806 311906 578830
rect 305938 572886 305962 578806
rect 307807 572886 310694 576661
rect 311882 572886 311906 578806
rect 305938 572862 311906 572886
rect 305298 572383 305618 572787
rect 298994 572284 304962 572308
rect 298994 566364 299018 572284
rect 300301 566364 303188 572284
rect 304938 566364 304962 572284
rect 298994 566340 304962 566364
rect 298354 565861 298674 566265
rect 292050 565762 298018 565786
rect 292050 559842 292074 565762
rect 293516 559842 296403 565762
rect 297994 559842 298018 565762
rect 292050 559818 298018 559842
rect 291410 559541 291730 559743
rect 259666 540435 259862 555640
rect 275226 540435 275332 555640
rect 229967 540409 229991 540415
rect 199671 540385 229991 540409
rect 128823 540159 131710 540383
rect 135608 540308 138495 540383
rect 149754 540308 152641 540383
rect 156683 540308 159570 540383
rect 100463 417422 101051 432558
rect 116402 417422 116619 432558
rect 100463 151638 116619 417422
rect 259666 378759 275332 540435
rect 293516 555337 296403 559818
rect 298354 559743 298396 565861
rect 298632 559743 298674 565861
rect 300301 565786 303188 566340
rect 305298 566265 305340 572383
rect 305576 566265 305618 572383
rect 307807 572308 310694 572862
rect 312242 572787 312284 578905
rect 312520 572787 312562 578905
rect 319186 578905 319506 583473
rect 312882 578806 318850 578830
rect 312882 572886 312906 578806
rect 314447 572886 317334 576733
rect 318826 572886 318850 578806
rect 312882 572862 318850 572886
rect 312242 572383 312562 572787
rect 305938 572284 311906 572308
rect 305938 566364 305962 572284
rect 307807 566364 310694 572284
rect 311882 566364 311906 572284
rect 305938 566340 311906 566364
rect 305298 565861 305618 566265
rect 298994 565762 304962 565786
rect 298994 559842 299018 565762
rect 300301 559842 303188 565762
rect 304938 559842 304962 565762
rect 298994 559818 304962 559842
rect 298354 559541 298674 559743
rect 300301 555337 303188 559818
rect 305298 559743 305340 565861
rect 305576 559743 305618 565861
rect 307807 565786 310694 566340
rect 312242 566265 312284 572383
rect 312520 566265 312562 572383
rect 314447 572308 317334 572862
rect 319186 572787 319228 578905
rect 319464 572787 319506 578905
rect 319826 578806 325794 578830
rect 319826 572886 319850 578806
rect 321376 572886 324263 576444
rect 325770 572886 325794 578806
rect 319826 572862 325794 572886
rect 319186 572383 319506 572787
rect 312882 572284 318850 572308
rect 312882 566364 312906 572284
rect 314447 566364 317334 572284
rect 318826 566364 318850 572284
rect 312882 566340 318850 566364
rect 312242 565861 312562 566265
rect 305938 565762 311906 565786
rect 305938 559842 305962 565762
rect 307807 559842 310694 565762
rect 311882 559842 311906 565762
rect 305938 559818 311906 559842
rect 305298 559541 305618 559743
rect 307807 555337 310694 559818
rect 312242 559743 312284 565861
rect 312520 559743 312562 565861
rect 314447 565786 317334 566340
rect 319186 566265 319228 572383
rect 319464 566265 319506 572383
rect 321376 572308 324263 572862
rect 319826 572284 325794 572308
rect 319826 566364 319850 572284
rect 321376 566364 324263 572284
rect 325770 566364 325794 572284
rect 319826 566340 325794 566364
rect 319186 565861 319506 566265
rect 312882 565762 318850 565786
rect 312882 559842 312906 565762
rect 314447 559842 317334 565762
rect 318826 559842 318850 565762
rect 312882 559818 318850 559842
rect 312242 559541 312562 559743
rect 314447 555337 317334 559818
rect 319186 559743 319228 565861
rect 319464 559743 319506 565861
rect 321376 565786 324263 566340
rect 319826 565762 325794 565786
rect 319826 559842 319850 565762
rect 321376 559842 324263 565762
rect 325770 559842 325794 565762
rect 319826 559818 325794 559842
rect 319186 559541 319506 559743
rect 321376 555337 324263 559818
rect 293516 555313 324263 555337
rect 293516 540369 293791 555313
rect 324068 540392 324263 555313
rect 324068 540369 324092 540392
rect 293516 540345 324092 540369
rect 293516 540198 296403 540345
rect 314447 540295 317334 540345
rect 259666 363295 259965 378759
rect 275183 363295 275332 378759
rect 259666 240427 275332 363295
rect 259666 225941 259755 240427
rect 259731 225260 259755 225941
rect 275011 225941 275332 240427
rect 338385 432559 354541 583865
rect 380930 583555 381126 598681
rect 411023 583555 411047 599184
rect 380930 583531 411047 583555
rect 380930 579563 383133 583531
rect 380930 579361 383208 579563
rect 380930 573243 383133 579361
rect 383166 573243 383208 579361
rect 389832 579361 390152 583531
rect 383528 579262 389496 579286
rect 383528 573342 383552 579262
rect 384994 573342 387881 577261
rect 389472 573342 389496 579262
rect 383528 573318 389496 573342
rect 380930 572839 383208 573243
rect 380930 566721 383133 572839
rect 383166 566721 383208 572839
rect 384994 572764 387881 573318
rect 389832 573243 389874 579361
rect 390110 573243 390152 579361
rect 396776 579361 397096 583531
rect 390472 579262 396440 579286
rect 390472 573342 390496 579262
rect 391779 573342 394666 577045
rect 396416 573342 396440 579262
rect 390472 573318 396440 573342
rect 389832 572839 390152 573243
rect 383528 572740 389496 572764
rect 383528 566820 383552 572740
rect 384994 566820 387881 572740
rect 389472 566820 389496 572740
rect 383528 566796 389496 566820
rect 380930 566317 383208 566721
rect 380930 560498 383133 566317
rect 382888 560199 382930 560498
rect 383166 560199 383208 566317
rect 384994 566242 387881 566796
rect 389832 566721 389874 572839
rect 390110 566721 390152 572839
rect 391779 572764 394666 573318
rect 396776 573243 396818 579361
rect 397054 573243 397096 579361
rect 403720 579361 404040 583531
rect 397416 579262 403384 579286
rect 397416 573342 397440 579262
rect 399285 573342 402172 577117
rect 403360 573342 403384 579262
rect 397416 573318 403384 573342
rect 396776 572839 397096 573243
rect 390472 572740 396440 572764
rect 390472 566820 390496 572740
rect 391779 566820 394666 572740
rect 396416 566820 396440 572740
rect 390472 566796 396440 566820
rect 389832 566317 390152 566721
rect 383528 566218 389496 566242
rect 383528 560298 383552 566218
rect 384994 560298 387881 566218
rect 389472 560298 389496 566218
rect 383528 560274 389496 560298
rect 382888 559997 383208 560199
rect 384994 555612 387881 560274
rect 389832 560199 389874 566317
rect 390110 560199 390152 566317
rect 391779 566242 394666 566796
rect 396776 566721 396818 572839
rect 397054 566721 397096 572839
rect 399285 572764 402172 573318
rect 403720 573243 403762 579361
rect 403998 573243 404040 579361
rect 410664 579361 410984 583531
rect 404360 579262 410328 579286
rect 404360 573342 404384 579262
rect 405925 573342 408812 577189
rect 410304 573342 410328 579262
rect 404360 573318 410328 573342
rect 403720 572839 404040 573243
rect 397416 572740 403384 572764
rect 397416 566820 397440 572740
rect 399285 566820 402172 572740
rect 403360 566820 403384 572740
rect 397416 566796 403384 566820
rect 396776 566317 397096 566721
rect 390472 566218 396440 566242
rect 390472 560298 390496 566218
rect 391779 560298 394666 566218
rect 396416 560298 396440 566218
rect 390472 560274 396440 560298
rect 389832 559997 390152 560199
rect 391779 555612 394666 560274
rect 396776 560199 396818 566317
rect 397054 560199 397096 566317
rect 399285 566242 402172 566796
rect 403720 566721 403762 572839
rect 403998 566721 404040 572839
rect 405925 572764 408812 573318
rect 410664 573243 410706 579361
rect 410942 573243 410984 579361
rect 411304 579262 417272 579286
rect 411304 573342 411328 579262
rect 412854 573342 415741 576900
rect 417248 573342 417272 579262
rect 411304 573318 417272 573342
rect 410664 572839 410984 573243
rect 404360 572740 410328 572764
rect 404360 566820 404384 572740
rect 405925 566820 408812 572740
rect 410304 566820 410328 572740
rect 404360 566796 410328 566820
rect 403720 566317 404040 566721
rect 397416 566218 403384 566242
rect 397416 560298 397440 566218
rect 399285 560298 402172 566218
rect 403360 560298 403384 566218
rect 397416 560274 403384 560298
rect 396776 559997 397096 560199
rect 399285 555612 402172 560274
rect 403720 560199 403762 566317
rect 403998 560199 404040 566317
rect 405925 566242 408812 566796
rect 410664 566721 410706 572839
rect 410942 566721 410984 572839
rect 412854 572764 415741 573318
rect 411304 572740 417272 572764
rect 411304 566820 411328 572740
rect 412854 566820 415741 572740
rect 417248 566820 417272 572740
rect 411304 566796 417272 566820
rect 410664 566317 410984 566721
rect 404360 566218 410328 566242
rect 404360 560298 404384 566218
rect 405925 560298 408812 566218
rect 410304 560298 410328 566218
rect 404360 560274 410328 560298
rect 403720 559997 404040 560199
rect 405925 555612 408812 560274
rect 410664 560199 410706 566317
rect 410942 560199 410984 566317
rect 412854 566242 415741 566796
rect 411304 566218 417272 566242
rect 411304 560298 411328 566218
rect 412854 560298 415741 566218
rect 417248 560298 417272 566218
rect 411304 560274 417272 560298
rect 410664 559997 410984 560199
rect 412854 555612 415741 560274
rect 384994 555588 415741 555612
rect 384994 540644 385148 555588
rect 415425 540644 415741 555588
rect 384994 540633 415741 540644
rect 385124 540620 415741 540633
rect 391779 540524 394666 540620
rect 412854 540415 415741 540620
rect 451976 555601 467642 673047
rect 510306 599189 525839 696878
rect 487908 599165 525839 599189
rect 487908 598849 487932 599165
rect 487426 583536 487932 598849
rect 525630 583536 525839 599165
rect 546152 598800 561241 598824
rect 546152 598734 546176 598800
rect 487426 583512 525839 583536
rect 487426 580018 489629 583512
rect 487426 579816 489704 580018
rect 487426 573698 489629 579816
rect 489662 573698 489704 579816
rect 496328 579816 496648 583512
rect 490024 579717 495992 579741
rect 490024 573797 490048 579717
rect 491490 573797 494377 577716
rect 495968 573797 495992 579717
rect 490024 573773 495992 573797
rect 487426 573294 489704 573698
rect 487426 567176 489629 573294
rect 489662 567176 489704 573294
rect 491490 573219 494377 573773
rect 496328 573698 496370 579816
rect 496606 573698 496648 579816
rect 503272 579816 503592 583512
rect 510173 583472 525839 583512
rect 545384 584066 546176 598734
rect 561217 598734 561241 598800
rect 561217 584066 561540 598734
rect 496968 579717 502936 579741
rect 496968 573797 496992 579717
rect 498275 573797 501162 577500
rect 502912 573797 502936 579717
rect 496968 573773 502936 573797
rect 496328 573294 496648 573698
rect 490024 573195 495992 573219
rect 490024 567275 490048 573195
rect 491490 567275 494377 573195
rect 495968 567275 495992 573195
rect 490024 567251 495992 567275
rect 487426 566772 489704 567176
rect 487426 560953 489629 566772
rect 489384 560654 489426 560953
rect 489662 560654 489704 566772
rect 491490 566697 494377 567251
rect 496328 567176 496370 573294
rect 496606 567176 496648 573294
rect 498275 573219 501162 573773
rect 503272 573698 503314 579816
rect 503550 573698 503592 579816
rect 510216 579816 510536 583472
rect 503912 579717 509880 579741
rect 503912 573797 503936 579717
rect 505781 573797 508668 577572
rect 509856 573797 509880 579717
rect 503912 573773 509880 573797
rect 503272 573294 503592 573698
rect 496968 573195 502936 573219
rect 496968 567275 496992 573195
rect 498275 567275 501162 573195
rect 502912 567275 502936 573195
rect 496968 567251 502936 567275
rect 496328 566772 496648 567176
rect 490024 566673 495992 566697
rect 490024 560753 490048 566673
rect 491490 560753 494377 566673
rect 495968 560753 495992 566673
rect 490024 560729 495992 560753
rect 489384 560452 489704 560654
rect 338385 417742 338894 432559
rect 354227 417742 354541 432559
rect 275011 225260 275035 225941
rect 259731 225236 275035 225260
rect 100463 136586 100582 151638
rect 116556 136586 116619 151638
rect 338385 151653 354541 417742
rect 451976 540149 452164 555601
rect 467493 540149 467642 555601
rect 491490 555373 494377 560729
rect 496328 560654 496370 566772
rect 496606 560654 496648 566772
rect 498275 566697 501162 567251
rect 503272 567176 503314 573294
rect 503550 567176 503592 573294
rect 505781 573219 508668 573773
rect 510216 573698 510258 579816
rect 510494 573698 510536 579816
rect 517160 579816 517480 583472
rect 510856 579717 516824 579741
rect 510856 573797 510880 579717
rect 512421 573797 515308 577644
rect 516800 573797 516824 579717
rect 510856 573773 516824 573797
rect 510216 573294 510536 573698
rect 503912 573195 509880 573219
rect 503912 567275 503936 573195
rect 505781 567275 508668 573195
rect 509856 567275 509880 573195
rect 503912 567251 509880 567275
rect 503272 566772 503592 567176
rect 496968 566673 502936 566697
rect 496968 560753 496992 566673
rect 498275 560753 501162 566673
rect 502912 560753 502936 566673
rect 496968 560729 502936 560753
rect 496328 560452 496648 560654
rect 498275 555373 501162 560729
rect 503272 560654 503314 566772
rect 503550 560654 503592 566772
rect 505781 566697 508668 567251
rect 510216 567176 510258 573294
rect 510494 567176 510536 573294
rect 512421 573219 515308 573773
rect 517160 573698 517202 579816
rect 517438 573698 517480 579816
rect 517800 579717 523768 579741
rect 517800 573797 517824 579717
rect 519350 573797 522237 577355
rect 523744 573797 523768 579717
rect 517800 573773 523768 573797
rect 517160 573294 517480 573698
rect 510856 573195 516824 573219
rect 510856 567275 510880 573195
rect 512421 567275 515308 573195
rect 516800 567275 516824 573195
rect 510856 567251 516824 567275
rect 510216 566772 510536 567176
rect 503912 566673 509880 566697
rect 503912 560753 503936 566673
rect 505781 560753 508668 566673
rect 509856 560753 509880 566673
rect 503912 560729 509880 560753
rect 503272 560452 503592 560654
rect 505781 555373 508668 560729
rect 510216 560654 510258 566772
rect 510494 560654 510536 566772
rect 512421 566697 515308 567251
rect 517160 567176 517202 573294
rect 517438 567176 517480 573294
rect 519350 573219 522237 573773
rect 517800 573195 523768 573219
rect 517800 567275 517824 573195
rect 519350 567275 522237 573195
rect 523744 567275 523768 573195
rect 517800 567251 523768 567275
rect 517160 566772 517480 567176
rect 510856 566673 516824 566697
rect 510856 560753 510880 566673
rect 512421 560753 515308 566673
rect 516800 560753 516824 566673
rect 510856 560729 516824 560753
rect 510216 560452 510536 560654
rect 512421 555373 515308 560729
rect 517160 560654 517202 566772
rect 517438 560654 517480 566772
rect 519350 566697 522237 567251
rect 517800 566673 523768 566697
rect 517800 560753 517824 566673
rect 519350 560753 522237 566673
rect 523744 560753 523768 566673
rect 517800 560729 523768 560753
rect 517160 560452 517480 560654
rect 519350 555373 522237 560729
rect 491289 555349 522237 555373
rect 491289 540466 491313 555349
rect 521955 540466 522237 555349
rect 491289 540442 522237 540466
rect 519350 540149 522237 540442
rect 451976 378918 467642 540149
rect 451976 363464 452093 378918
rect 467213 363464 467642 378918
rect 451976 240355 467642 363464
rect 451976 227015 452031 240355
rect 452007 225376 452031 227015
rect 467535 227015 467642 240355
rect 545384 432093 561540 584066
rect 545384 417276 545705 432093
rect 561038 417276 561540 432093
rect 467535 225376 467559 227015
rect 452007 225352 467559 225376
rect 338385 136722 338641 151653
rect 100463 136311 116619 136586
rect 338617 136461 338641 136722
rect 354383 136722 354541 151653
rect 545384 151702 561540 417276
rect 545384 137728 545482 151702
rect 354383 136461 354407 136722
rect 545458 136619 545482 137728
rect 561448 137728 561540 151702
rect 561448 136619 561472 137728
rect 545458 136595 561472 136619
rect 338617 136437 354407 136461
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use mimcap_decoup_1x5  mimcap_decoup_1x5_0
array 0 0 34500 0 2 6522
timestamp 1624376995
transform 1 0 38481 0 1 560871
box 0 -159 34500 6363
use top_pll_v1  top_pll_v1_0
timestamp 1624402156
transform 1 0 14782 0 1 657248
box -642 -33679 50180 2860
use sky130_fd_pr__cap_mim_m3_2_2Y8F6P  sky130_fd_pr__cap_mim_m3_2_2Y8F6P_0
array 0 0 6724 0 8 6522
timestamp 1624129585
transform 1 0 74005 0 1 616157
box -3351 -3261 3373 3261
use top_pll_v2 *top_pll_v2_0
timestamp 1624402156
transform -1 0 133068 0 1 657248
box -642 -33679 50180 2860
use mimcap_decoup_1x5  mimcap_decoup_1x5_1
array 0 0 34500 0 2 6522
timestamp 1624376995
transform 1 0 126717 0 1 559996
box 0 -159 34500 6363
use sky130_fd_pr__cap_mim_m3_2_2Y8F6P  sky130_fd_pr__cap_mim_m3_2_2Y8F6P_1
array 0 0 6724 0 8 6522
timestamp 1624129585
transform 1 0 144463 0 1 616442
box -3351 -3261 3373 3261
use top_pll_v1 *top_pll_v1_1
timestamp 1624402156
transform -1 0 206380 0 1 656706
box -642 -33679 50180 2860
use sky130_fd_pr__cap_mim_m3_2_2Y8F6P  sky130_fd_pr__cap_mim_m3_2_2Y8F6P_2
array 0 0 6724 0 6 6522
timestamp 1624129585
transform 1 0 220679 0 1 616773
box -3351 -3261 3373 3261
use mimcap_decoup_1x5  mimcap_decoup_1x5_2
array 0 0 34500 0 2 6522
timestamp 1624376995
transform 1 0 197202 0 1 560156
box 0 -159 34500 6363
use bias  bias_0
timestamp 1624049879
transform 1 0 202834 0 -1 687483
box -54 -412 44317 2238
use mimcap_decoup_1x5  mimcap_decoup_1x5_6
array 0 0 34500 0 1 6522
timestamp 1624376995
transform -1 0 345445 0 1 602155
box 0 -159 34500 6363
use mimcap_decoup_1x5  mimcap_decoup_1x5_3
array 0 0 34500 0 2 6522
timestamp 1624376995
transform 1 0 291410 0 1 559700
box 0 -159 34500 6363
use res_amp_top  res_amp_top_0 ~/caravel_analog_fulgor/mag/afernandez_residue_amplifier
timestamp 1624402156
transform 1 0 349695 0 1 630386
box -5005 -972 31038 12726
use mimcap_decoup_1x5  mimcap_decoup_1x5_4
array 0 0 34500 0 2 6522
timestamp 1624376995
transform 1 0 382888 0 1 560156
box 0 -159 34500 6363
use mimcap_decoup_1x5  mimcap_decoup_1x5_5
array 0 0 34500 0 2 6522
timestamp 1624376995
transform 1 0 489384 0 1 560611
box 0 -159 34500 6363
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s -800 559442 860 564242 0 FreeSans 1120 180 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
