magic
tech sky130A
magscale 1 2
timestamp 1624396964
<< nwell >>
rect 0 2846 20536 2860
rect 0 2838 6183 2846
rect 0 2608 3909 2838
rect 3790 2062 3909 2608
rect 6063 2012 6183 2838
rect 13905 2752 20536 2846
rect 13905 1955 14025 2752
rect 18329 1955 20536 2752
rect 18510 1923 20536 1955
rect 20472 1290 20536 1923
rect 49317 1290 50180 2860
rect -3 -230 3909 546
rect -3 -350 6063 -230
rect 955 -370 2001 -350
<< pwell >>
rect 3790 706 3909 2062
rect 2872 546 3909 706
rect 13905 784 14901 854
rect 18329 784 18510 1215
rect 20472 1190 20593 1290
rect 20456 1176 20593 1190
rect 13905 653 18510 784
rect 19367 653 20225 754
rect 20472 653 20593 1176
rect 13905 223 20593 653
rect 13905 181 20796 223
rect 27347 181 46785 1226
rect 49317 769 50180 1290
rect 49319 181 50180 769
rect 13905 -238 50180 181
rect 19278 -3693 50180 -238
rect 19278 -3827 49370 -3693
rect 20572 -4375 49370 -3827
<< psubdiff >>
rect 20575 24 20599 114
rect 49259 24 49283 114
rect 48569 -453 50169 -429
rect 13461 -1919 13485 -1831
rect 14493 -1919 14517 -1831
rect 48569 -4056 50169 -4032
<< nsubdiff >>
rect 43 -212 67 -124
rect 416 -212 440 -124
rect 1252 -220 1276 -132
rect 1625 -220 1649 -132
rect 2420 -214 2446 -126
rect 2795 -214 2819 -126
<< psubdiffcont >>
rect 20599 24 49259 114
rect 13485 -1919 14493 -1831
rect 48569 -4032 50169 -453
<< nsubdiffcont >>
rect 67 -212 416 -124
rect 1276 -220 1625 -132
rect 2446 -214 2795 -126
<< poly >>
rect 10374 2156 10680 2179
rect 10374 2078 10395 2156
rect 10657 2078 10680 2156
rect 10374 2055 10680 2078
rect 10354 385 10697 405
rect 10354 280 10372 385
rect 10671 280 10697 385
rect 10354 269 10697 280
<< polycont >>
rect 9420 2020 9699 2114
rect 10395 2078 10657 2156
rect 9434 325 9696 449
rect 10372 280 10671 385
<< locali >>
rect 20583 24 20599 114
rect 49259 24 49275 114
rect 48569 -453 50169 -437
rect 48569 -4048 50169 -4032
<< viali >>
rect 10374 2156 10680 2179
rect 9399 2114 9723 2134
rect 9399 2020 9420 2114
rect 9420 2020 9699 2114
rect 9699 2020 9723 2114
rect 10374 2078 10395 2156
rect 10395 2078 10657 2156
rect 10657 2078 10680 2156
rect 10374 2055 10680 2078
rect 9399 1999 9723 2020
rect 9405 449 9723 468
rect 9405 325 9434 449
rect 9434 325 9696 449
rect 9696 325 9723 449
rect 9405 306 9723 325
rect 10354 385 10697 405
rect 10354 280 10372 385
rect 10372 280 10671 385
rect 10671 280 10697 385
rect 10354 269 10697 280
rect 20599 24 49259 114
rect 22 -124 2852 -112
rect 22 -212 67 -124
rect 67 -212 416 -124
rect 416 -126 2852 -124
rect 416 -132 2446 -126
rect 416 -212 1276 -132
rect 22 -220 1276 -212
rect 1276 -220 1625 -132
rect 1625 -214 2446 -132
rect 2446 -214 2795 -126
rect 2795 -214 2852 -126
rect 1625 -220 2852 -214
rect 22 -232 2852 -220
rect 13416 -1831 14548 -1810
rect 13416 -1919 13485 -1831
rect 13485 -1919 14493 -1831
rect 14493 -1919 14548 -1831
rect 13416 -1931 14548 -1919
rect 48569 -4032 50169 -453
<< metal1 >>
rect 0 2824 20536 2830
rect 0 2816 20548 2824
rect 0 2808 6183 2816
rect 0 2674 6294 2808
rect 13869 2687 20548 2816
rect 13869 2674 20472 2687
rect 0 2578 3504 2674
rect 3150 2150 3504 2578
rect 5909 2095 6099 2096
rect 4963 2090 5581 2095
rect 3909 2034 3919 2090
rect 4143 2034 4153 2090
rect 4963 2034 5180 2090
rect 5404 2034 5581 2090
rect 4963 2029 5581 2034
rect 5873 2091 6099 2095
rect 5873 2035 5955 2091
rect 6089 2035 6099 2091
rect 5873 2030 6099 2035
rect 5873 2029 6063 2030
rect 0 1956 210 2022
rect 8859 2012 8963 2633
rect 13835 2624 20472 2674
rect 13835 2617 14025 2624
rect 10362 2179 10692 2185
rect 9387 2134 9735 2140
rect 9387 1999 9399 2134
rect 9723 1999 9735 2134
rect 10362 2055 10374 2179
rect 10680 2055 10692 2179
rect 11133 2158 11217 2499
rect 10362 2049 10692 2055
rect 9387 1993 9735 1999
rect 18308 1990 20472 2624
rect 18329 1985 20472 1990
rect 18510 1880 20472 1985
rect 18510 1879 19087 1880
rect 18863 1841 19087 1879
rect 18863 1823 19020 1841
rect 3857 1234 3909 1468
rect 6052 1268 6259 1468
rect 3857 870 3976 1234
rect 3790 830 3976 870
rect 3585 776 3976 830
rect 3790 736 3976 776
rect 6183 830 6259 1268
rect 18510 1190 18520 1242
rect 18728 1190 18738 1242
rect 18878 1176 19279 1256
rect 19577 1172 19587 1256
rect 19999 1172 20009 1256
rect 20308 1250 20318 1253
rect 20305 1172 20318 1250
rect 20308 1169 20318 1172
rect 20560 1241 20570 1253
rect 20560 1182 20839 1241
rect 20560 1169 20570 1182
rect 48286 1072 49317 1356
rect -619 518 -609 715
rect -513 652 -503 715
rect 6183 695 6219 830
rect 18329 723 18510 783
rect 18326 715 19398 723
rect 18326 712 19370 715
rect -513 586 210 652
rect -513 518 -503 586
rect 5003 574 5581 579
rect 3909 518 3919 574
rect 4143 518 4153 574
rect 5003 518 5180 574
rect 5404 518 5581 574
rect 5003 513 5581 518
rect 5873 574 6063 579
rect 5873 518 5919 574
rect 6053 518 6063 574
rect 5873 513 6063 518
rect 9393 468 9735 474
rect 6405 392 8963 408
rect 6403 320 8963 392
rect 6405 304 8963 320
rect 9393 306 9405 468
rect 9723 306 9735 468
rect 9393 300 9735 306
rect 10342 405 10709 411
rect 10342 269 10354 405
rect 10697 269 10709 405
rect 10342 263 10709 269
rect -1 -106 499 93
rect 1102 19 1997 124
rect 11118 80 11244 311
rect 1194 -106 1694 19
rect 2372 -106 2872 55
rect 18326 -66 19612 712
rect 20472 677 20536 788
rect 20443 244 20536 677
rect 24126 244 24570 245
rect 48566 244 49046 267
rect 20443 114 49287 244
rect 20443 24 20599 114
rect 49259 24 49287 114
rect 20443 18 49287 24
rect -1 -112 2872 -106
rect -1 -232 22 -112
rect 2852 -232 2872 -112
rect -1 -238 2872 -232
rect -1 -407 499 -238
rect 1194 -370 1694 -238
rect 1102 -514 1997 -370
rect 2372 -445 2872 -238
rect 3909 -380 6063 -200
rect 13905 -208 19612 -66
rect -627 -1095 -617 -882
rect -505 -1095 -495 -882
rect 6175 -1110 6996 -1051
rect 13787 -1223 13797 -1056
rect 13962 -1092 13972 -1056
rect 13962 -1170 13973 -1092
rect 14281 -1166 14682 -1086
rect 14819 -1154 15043 -1098
rect 13962 -1223 13972 -1170
rect 13580 -1706 13842 -1507
rect 13580 -1725 14356 -1706
rect 19367 -1720 19612 -208
rect 48566 -441 49046 18
rect 13288 -1896 13289 -1731
rect 13768 -1804 14356 -1725
rect 13404 -1810 14560 -1804
rect 13404 -1931 13416 -1810
rect 14548 -1931 14560 -1810
rect 13404 -1937 14560 -1931
rect 13768 -2069 14356 -1937
rect 19278 -1964 19612 -1720
rect 48563 -453 50175 -441
rect 13768 -2215 13842 -2069
rect 10227 -2717 10598 -2658
rect 13760 -2695 13770 -2498
rect 13951 -2599 13961 -2498
rect 13951 -2677 13973 -2599
rect 13951 -2695 13961 -2677
rect 14281 -2683 14682 -2603
rect 14816 -2673 15040 -2617
rect 48563 -4032 48569 -453
rect 50169 -4032 50175 -453
rect 48563 -5101 50175 -4032
<< via1 >>
rect 3919 2034 4143 2090
rect 5180 2034 5404 2090
rect 5955 2035 6089 2091
rect 9420 2020 9699 2114
rect 10395 2078 10657 2156
rect 18520 1190 18728 1242
rect 19587 1172 19999 1256
rect 20318 1169 20560 1253
rect -609 518 -513 715
rect 3919 518 4143 574
rect 5180 518 5404 574
rect 5919 518 6053 574
rect 9434 325 9696 449
rect 10372 280 10671 385
rect -617 -1095 -505 -882
rect 13797 -1223 13962 -1056
rect 13770 -2695 13951 -2498
<< metal2 >>
rect 10395 2156 10657 2166
rect 9420 2114 9699 2124
rect 3919 2090 4143 2100
rect 3919 2024 4143 2034
rect 5180 2090 5404 2100
rect 5180 2024 5404 2034
rect 5955 2091 6089 2101
rect 5955 2025 6089 2035
rect 10395 2068 10657 2078
rect 3988 1928 4074 2024
rect 9420 2010 9699 2020
rect 3738 1876 4074 1928
rect 5955 1831 9647 1854
rect 5955 1812 9499 1831
rect 6089 1775 9499 1812
rect 9633 1775 9647 1831
rect 6089 1756 9647 1775
rect 2159 858 2211 1750
rect 5955 1746 9647 1756
rect 5232 1611 10645 1637
rect 5232 1555 5245 1611
rect 5469 1609 10645 1611
rect 5469 1555 10410 1609
rect 5232 1553 10410 1555
rect 10634 1553 10645 1609
rect 5232 1529 10645 1553
rect 19587 1256 19999 1266
rect 18520 1242 18728 1252
rect 18091 1190 18520 1241
rect 18091 1189 18728 1190
rect 18520 1180 18728 1189
rect 19587 1162 19999 1172
rect 20318 1253 20560 1263
rect 20318 1159 20560 1169
rect 5232 1055 10645 1079
rect 5232 1053 10410 1055
rect 5232 997 5245 1053
rect 5469 999 10410 1053
rect 10634 999 10645 1055
rect 5469 997 10645 999
rect 5232 971 10645 997
rect 13187 980 13690 990
rect 5919 853 9631 863
rect 6053 797 9497 853
rect 5919 755 9631 797
rect 3988 732 4074 733
rect -609 715 -513 725
rect 3685 680 4074 732
rect 3988 584 4074 680
rect -609 508 -513 518
rect 3919 574 4143 584
rect 3919 508 4143 518
rect 5180 574 5404 584
rect 5180 508 5404 518
rect 5919 574 6053 584
rect 5919 508 6053 518
rect 9434 449 9696 459
rect 9434 315 9696 325
rect 10372 385 10671 395
rect 13187 381 13690 391
rect 10372 270 10671 280
rect 13764 206 14377 369
rect 14214 25 14377 206
rect -617 -882 -505 -872
rect -279 -954 161 -878
rect -617 -1105 -505 -1095
rect 13797 -1056 13962 -1046
rect -405 -1940 -319 -1188
rect 13797 -1233 13962 -1223
rect 9937 -2546 10013 -1824
rect 13770 -2498 13951 -2488
rect 13770 -2705 13951 -2695
<< via2 >>
rect 5180 2034 5404 2090
rect 5955 2035 6089 2091
rect 9491 2043 9625 2099
rect 10412 2078 10636 2134
rect 5955 1756 6089 1812
rect 9499 1775 9633 1831
rect 5245 1555 5469 1611
rect 10410 1553 10634 1609
rect 19587 1172 19999 1256
rect 5245 997 5469 1053
rect 10410 999 10634 1055
rect 5919 797 6053 853
rect 9497 797 9631 853
rect -609 518 -513 715
rect 5180 518 5404 574
rect 5919 518 6053 574
rect 9497 359 9631 415
rect 13187 391 13690 980
rect 10412 306 10636 362
rect -617 -1095 -505 -882
rect 13797 -1223 13962 -1056
rect 13770 -2695 13951 -2498
<< metal3 >>
rect 10402 2134 10646 2139
rect 9470 2099 9672 2114
rect 5170 2090 5414 2095
rect 5170 2034 5180 2090
rect 5404 2034 5414 2090
rect 5170 2029 5414 2034
rect 5945 2091 6099 2096
rect 5945 2035 5955 2091
rect 6089 2035 6099 2091
rect 5945 2030 6099 2035
rect 9470 2043 9491 2099
rect 9625 2043 9672 2099
rect 10402 2078 10412 2134
rect 10636 2078 10646 2134
rect 10402 2073 10646 2078
rect 9470 2034 9672 2043
rect 5262 1616 5322 2029
rect 5992 1817 6052 2030
rect 9525 1836 9585 2034
rect 9489 1831 9643 1836
rect 5945 1812 6099 1817
rect 5945 1756 5955 1812
rect 6089 1756 6099 1812
rect 9489 1775 9499 1831
rect 9633 1775 9643 1831
rect 9489 1770 9643 1775
rect 9525 1769 9585 1770
rect 5945 1751 6099 1756
rect 5992 1742 6052 1751
rect 5235 1611 5479 1616
rect 10494 1614 10554 2073
rect 5235 1555 5245 1611
rect 5469 1555 5479 1611
rect 5235 1550 5479 1555
rect 10400 1609 10644 1614
rect 10400 1553 10410 1609
rect 10634 1553 10644 1609
rect 10400 1548 10644 1553
rect 19577 1256 20009 1261
rect 19577 1172 19587 1256
rect 19999 1172 20009 1256
rect 19577 1167 20009 1172
rect 5235 1053 5479 1058
rect 5235 997 5245 1053
rect 5469 997 5479 1053
rect 5235 992 5479 997
rect 10400 1055 10644 1060
rect 10400 999 10410 1055
rect 10634 999 10644 1055
rect 10400 994 10644 999
rect -627 715 -495 725
rect -627 518 -609 715
rect -513 518 -495 715
rect 5262 579 5322 992
rect 5956 858 6016 867
rect 5909 853 6063 858
rect 5909 797 5919 853
rect 6053 797 6063 853
rect 5909 792 6063 797
rect 9487 853 9641 858
rect 9487 797 9497 853
rect 9631 797 9641 853
rect 9487 792 9641 797
rect 5956 579 6016 792
rect -627 -882 -495 518
rect 5170 574 5414 579
rect 5170 518 5180 574
rect 5404 518 5414 574
rect 5170 513 5414 518
rect 5909 574 6063 579
rect 5909 518 5919 574
rect 6053 518 6063 574
rect 5909 513 6063 518
rect 9534 420 9594 792
rect 9487 415 9641 420
rect 9487 359 9497 415
rect 9631 359 9641 415
rect 10494 367 10554 994
rect 13177 980 13700 985
rect 13177 391 13187 980
rect 13690 391 13700 980
rect 13177 386 13700 391
rect 9487 354 9641 359
rect 10402 362 10646 367
rect 10402 306 10412 362
rect 10636 306 10646 362
rect 10402 301 10646 306
rect -627 -1095 -617 -882
rect -505 -1095 -495 -882
rect -627 -1100 -495 -1095
rect 13224 -3781 13580 386
rect 16756 -71 16812 -15
rect 13787 -1053 13972 -1051
rect 13785 -1259 13795 -1053
rect 13965 -1259 13975 -1053
rect 18944 -1835 19058 -1290
rect 18937 -1939 18947 -1835
rect 19055 -1939 19065 -1835
rect 19758 -1841 19952 1167
rect 19758 -1930 19773 -1841
rect 19940 -1930 19952 -1841
rect 13760 -2498 13961 -2493
rect 13760 -2695 13770 -2498
rect 13951 -2695 13961 -2498
rect 13760 -2700 13961 -2695
rect 18944 -2750 19058 -1939
rect 19758 -1964 19952 -1930
rect 13067 -4358 13077 -3781
rect 13764 -4358 13774 -3781
<< via3 >>
rect 13795 -1056 13965 -1053
rect 13795 -1223 13797 -1056
rect 13797 -1223 13962 -1056
rect 13962 -1223 13965 -1056
rect 13795 -1259 13965 -1223
rect 18947 -1939 19055 -1835
rect 19773 -1930 19940 -1841
rect 13770 -2695 13951 -2498
rect 13077 -4358 13764 -3781
<< metal4 >>
rect 638 -1053 13971 -1048
rect 638 -1259 13795 -1053
rect 13965 -1259 13971 -1053
rect 638 -1271 13971 -1259
rect 18944 -1835 19952 -1831
rect 18944 -1939 18947 -1835
rect 19055 -1841 19952 -1835
rect 19055 -1930 19773 -1841
rect 19940 -1930 19952 -1841
rect 19055 -1939 19952 -1930
rect 18944 -1943 19952 -1939
rect 638 -2498 13971 -2481
rect 638 -2695 13770 -2498
rect 13951 -2695 13971 -2498
rect 638 -2704 13971 -2695
rect 13076 -3781 13765 -3780
rect 13076 -4358 13077 -3781
rect 13764 -4358 13765 -3781
rect 13076 -4359 13765 -4358
rect 19686 -4493 43939 -3693
use loop_filter  loop_filter_0
timestamp 1624049879
transform 1 0 15820 0 1 -9473
box -16462 -24206 34360 5780
use charge_pump  charge_pump_0
timestamp 1624049879
transform 1 0 6183 0 1 -142
box 0 -96 7722 2988
use buffer_salida  buffer_salida_0
timestamp 1624049879
transform 1 0 20599 0 1 1292
box -63 -1119 28718 1568
use pfd_cp_interface  pfd_cp_interface_0
timestamp 1624049879
transform 1 0 3909 0 1 -230
box 0 0 2154 3068
use PFD  PFD_0
timestamp 1624049879
transform 1 0 0 0 1 1304
box 0 -1304 3790 1304
use ring_osc  ring_osc_0
timestamp 1624049879
transform 1 0 14447 0 1 -174
box -422 0 3882 2956
use ring_osc_buffer  ring_osc_buffer_0
timestamp 1624396964
transform 1 0 18509 0 1 653
box 0 0 1963 1270
use div_by_5  div_by_5_0
timestamp 1624396964
transform -1 0 13250 0 1 -3418
box -556 0 13892 3068
use div_by_2  div_by_2_0
timestamp 1624396964
transform -1 0 18034 0 -1 -350
box -1244 0 4228 3068
<< labels >>
rlabel metal2 2159 858 2211 1750 1 pfd_reset
rlabel metal1 0 1956 210 2022 1 in_ref
rlabel metal2 3988 1876 4074 2034 1 QA
rlabel metal2 3988 574 4074 733 1 QB
rlabel metal2 6053 755 9497 863 1 Down
rlabel metal2 5469 971 10410 1079 1 nDown
rlabel metal2 5469 1529 10410 1637 1 Up
rlabel metal2 6089 1746 9499 1854 1 nUp
rlabel metal1 8859 2012 8963 2633 1 biasp
rlabel metal1 11133 2158 11217 2499 1 pswitch
rlabel metal1 11118 80 11244 311 1 nswitch
rlabel metal2 13764 206 14377 369 1 vco_vctrl
rlabel metal3 16756 -71 16812 -15 1 vco_D0
rlabel metal2 18091 1189 18520 1241 1 vco_out
rlabel metal1 18878 1176 19279 1256 1 out_first_buffer
rlabel via1 19587 1172 19999 1256 1 out_to_div
rlabel metal1 14816 -2673 15040 -2617 1 out_div_2
rlabel metal1 14819 -1154 15043 -1098 1 n_out_div_2
rlabel metal1 14281 -1166 14682 -1086 1 n_out_buffer_div_2
rlabel metal1 14281 -2683 14682 -2603 1 out_buffer_div_2
rlabel metal1 13806 -2677 13973 -2599 1 out_by_2
rlabel metal1 13806 -1170 13973 -1092 1 n_out_by_2
rlabel metal2 -279 -954 161 -878 1 div_5_Q1_shift
rlabel metal3 -627 -882 -495 518 1 out_div_by_5
rlabel metal2 -405 -1940 -319 -1188 1 div_5_Q1
rlabel metal1 6175 -1110 6996 -1051 1 div_5_Q0
rlabel metal2 9937 -2546 10013 -1824 1 div_5_nQ0
rlabel metal1 10227 -2717 10598 -2658 1 div_5_nQ2
rlabel metal1 6405 304 8963 408 1 iref_cp
rlabel metal1 0 2578 3504 2816 1 vdd
rlabel metal1 18326 -208 19370 723 1 vss
rlabel metal4 19686 -4493 43939 -3693 1 lf_vc
rlabel metal1 20560 1182 20839 1241 1 out_to_buffer
rlabel metal1 48286 1072 49317 1356 1 out_to_pad
<< end >>
