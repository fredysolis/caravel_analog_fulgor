magic
tech sky130A
timestamp 1623247475
<< metal1 >>
rect 317 231 357 257
rect 383 231 423 257
rect 317 229 343 231
rect 277 177 303 217
rect 277 125 303 151
rect 277 73 303 99
rect 277 23 303 47
rect 397 229 423 231
rect 317 177 343 203
rect 317 125 343 151
rect 317 73 343 99
rect 317 37 343 47
rect 357 177 383 217
rect 357 125 383 151
rect 357 73 383 99
rect 357 23 383 47
rect 397 177 423 203
rect 397 125 423 151
rect 397 73 423 99
rect 397 37 423 47
rect 437 177 463 217
rect 437 125 463 151
rect 437 73 463 99
rect 437 23 463 47
rect 277 -3 317 23
rect 343 -3 397 23
rect 423 -3 463 23
<< via1 >>
rect 357 231 383 257
rect 277 151 303 177
rect 277 99 303 125
rect 277 47 303 73
rect 317 203 343 229
rect 317 151 343 177
rect 317 99 343 125
rect 317 47 343 73
rect 357 151 383 177
rect 357 99 383 125
rect 357 47 383 73
rect 397 203 423 229
rect 397 151 423 177
rect 397 99 423 125
rect 397 47 423 73
rect 437 151 463 177
rect 437 99 463 125
rect 437 47 463 73
rect 317 -3 343 23
rect 397 -3 423 23
<< metal2 >>
rect 317 231 357 257
rect 383 231 423 257
rect 317 229 343 231
rect 277 177 303 217
rect 277 125 303 151
rect 277 73 303 99
rect 277 23 303 47
rect 397 229 423 231
rect 317 177 343 203
rect 317 125 343 151
rect 317 73 343 99
rect 317 37 343 47
rect 357 177 383 217
rect 357 125 383 151
rect 357 73 383 99
rect 357 23 383 47
rect 397 177 423 203
rect 397 125 423 151
rect 397 73 423 99
rect 397 37 423 47
rect 437 177 463 217
rect 437 125 463 151
rect 437 73 463 99
rect 437 23 463 47
rect 277 -3 317 23
rect 343 -3 397 23
rect 423 -3 463 23
<< labels >>
rlabel via1 357 231 383 257 1 b
rlabel metal2 357 -3 383 23 1 t
<< end >>
