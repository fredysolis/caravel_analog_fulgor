magic
tech sky130A
magscale 1 2
timestamp 1622843784
<< pwell >>
rect -647 -360 647 360
<< nmos >>
rect -447 -150 -417 150
rect -351 -150 -321 150
rect -255 -150 -225 150
rect -159 -150 -129 150
rect -63 -150 -33 150
rect 33 -150 63 150
rect 129 -150 159 150
rect 225 -150 255 150
rect 321 -150 351 150
rect 417 -150 447 150
<< ndiff >>
rect -509 138 -447 150
rect -509 -138 -497 138
rect -463 -138 -447 138
rect -509 -150 -447 -138
rect -417 138 -351 150
rect -417 -138 -401 138
rect -367 -138 -351 138
rect -417 -150 -351 -138
rect -321 138 -255 150
rect -321 -138 -305 138
rect -271 -138 -255 138
rect -321 -150 -255 -138
rect -225 138 -159 150
rect -225 -138 -209 138
rect -175 -138 -159 138
rect -225 -150 -159 -138
rect -129 138 -63 150
rect -129 -138 -113 138
rect -79 -138 -63 138
rect -129 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 129 150
rect 63 -138 79 138
rect 113 -138 129 138
rect 63 -150 129 -138
rect 159 138 225 150
rect 159 -138 175 138
rect 209 -138 225 138
rect 159 -150 225 -138
rect 255 138 321 150
rect 255 -138 271 138
rect 305 -138 321 138
rect 255 -150 321 -138
rect 351 138 417 150
rect 351 -138 367 138
rect 401 -138 417 138
rect 351 -150 417 -138
rect 447 138 509 150
rect 447 -138 463 138
rect 497 -138 509 138
rect 447 -150 509 -138
<< ndiffc >>
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
<< psubdiff >>
rect -611 290 -515 324
rect 515 290 611 324
rect -611 228 -577 290
rect 577 228 611 290
rect -611 -290 -577 -228
rect 577 -290 611 -228
rect -611 -324 -515 -290
rect 515 -324 611 -290
<< psubdiffcont >>
rect -515 290 515 324
rect -611 -228 -577 228
rect 577 -228 611 228
rect -515 -324 515 -290
<< poly >>
rect -465 222 465 238
rect -465 188 -449 222
rect -415 188 -353 222
rect -319 188 -257 222
rect -223 188 -161 222
rect -127 188 -65 222
rect -31 188 31 222
rect 65 188 127 222
rect 161 188 223 222
rect 257 188 319 222
rect 353 188 415 222
rect 449 188 465 222
rect -465 172 465 188
rect -447 150 -417 172
rect -351 150 -321 172
rect -255 150 -225 172
rect -159 150 -129 172
rect -63 150 -33 172
rect 33 150 63 172
rect 129 150 159 172
rect 225 150 255 172
rect 321 150 351 172
rect 417 150 447 172
rect -447 -176 -417 -150
rect -351 -176 -321 -150
rect -255 -176 -225 -150
rect -159 -176 -129 -150
rect -63 -176 -33 -150
rect 33 -176 63 -150
rect 129 -176 159 -150
rect 225 -176 255 -150
rect 321 -176 351 -150
rect 417 -176 447 -150
<< polycont >>
rect -449 188 -415 222
rect -353 188 -319 222
rect -257 188 -223 222
rect -161 188 -127 222
rect -65 188 -31 222
rect 31 188 65 222
rect 127 188 161 222
rect 223 188 257 222
rect 319 188 353 222
rect 415 188 449 222
<< locali >>
rect -611 290 -515 324
rect 515 290 611 324
rect -611 228 -577 290
rect 577 228 611 290
rect -465 188 -449 222
rect -415 188 -353 222
rect -319 188 -257 222
rect -223 188 -161 222
rect -127 188 -65 222
rect -31 188 31 222
rect 65 188 127 222
rect 161 188 223 222
rect 257 188 319 222
rect 353 188 415 222
rect 449 188 465 222
rect -497 138 -463 154
rect -497 -154 -463 -138
rect -401 138 -367 154
rect -401 -154 -367 -138
rect -305 138 -271 154
rect -305 -154 -271 -138
rect -209 138 -175 154
rect -209 -154 -175 -138
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect 175 138 209 154
rect 175 -154 209 -138
rect 271 138 305 154
rect 271 -154 305 -138
rect 367 138 401 154
rect 367 -154 401 -138
rect 463 138 497 154
rect 463 -154 497 -138
rect -611 -290 -577 -228
rect 577 -290 611 -228
rect -611 -324 -515 -290
rect 515 -324 611 -290
<< viali >>
rect -449 188 -415 222
rect -353 188 -319 222
rect -257 188 -223 222
rect -161 188 -127 222
rect -65 188 -31 222
rect 31 188 65 222
rect 127 188 161 222
rect 223 188 257 222
rect 319 188 353 222
rect 415 188 449 222
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
<< metal1 >>
rect -464 222 464 231
rect -464 188 -449 222
rect -415 188 -353 222
rect -319 188 -257 222
rect -223 188 -161 222
rect -127 188 -65 222
rect -31 188 31 222
rect 65 188 127 222
rect 161 188 223 222
rect 257 188 319 222
rect 353 188 415 222
rect 449 188 464 222
rect -464 179 464 188
rect -503 138 -457 150
rect -503 -138 -497 138
rect -463 -138 -457 138
rect -503 -150 -457 -138
rect -407 138 -361 150
rect -407 -138 -401 138
rect -367 -138 -361 138
rect -407 -150 -361 -138
rect -311 138 -265 150
rect -311 -138 -305 138
rect -271 -138 -265 138
rect -311 -150 -265 -138
rect -215 138 -169 150
rect -215 -138 -209 138
rect -175 -138 -169 138
rect -215 -150 -169 -138
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -150 -73 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -150 119 -138
rect 169 138 215 150
rect 169 -138 175 138
rect 209 -138 215 138
rect 169 -150 215 -138
rect 265 138 311 150
rect 265 -138 271 138
rect 305 -138 311 138
rect 265 -150 311 -138
rect 361 138 407 150
rect 361 -138 367 138
rect 401 -138 407 138
rect 361 -150 407 -138
rect 457 138 503 150
rect 457 -138 463 138
rect 497 -138 503 138
rect 457 -150 503 -138
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -594 -307 594 307
string parameters w 1.5 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
