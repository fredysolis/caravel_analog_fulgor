magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect -359 -303 359 303
<< pmos >>
rect -159 -84 -129 84
rect -63 -84 -33 84
rect 33 -84 63 84
rect 129 -84 159 84
<< pdiff >>
rect -221 72 -159 84
rect -221 -72 -209 72
rect -175 -72 -159 72
rect -221 -84 -159 -72
rect -129 72 -63 84
rect -129 -72 -113 72
rect -79 -72 -63 72
rect -129 -84 -63 -72
rect -33 72 33 84
rect -33 -72 -17 72
rect 17 -72 33 72
rect -33 -84 33 -72
rect 63 72 129 84
rect 63 -72 79 72
rect 113 -72 129 72
rect 63 -84 129 -72
rect 159 72 221 84
rect 159 -72 175 72
rect 209 -72 221 72
rect 159 -84 221 -72
<< pdiffc >>
rect -209 -72 -175 72
rect -113 -72 -79 72
rect -17 -72 17 72
rect 79 -72 113 72
rect 175 -72 209 72
<< nsubdiff >>
rect -323 233 -227 267
rect 227 233 323 267
rect -323 171 -289 233
rect 289 171 323 233
rect -323 -233 -289 -171
rect 289 -233 323 -171
<< nsubdiffcont >>
rect -227 233 227 267
rect -323 -171 -289 171
rect 289 -171 323 171
<< poly >>
rect -159 84 -129 110
rect -63 84 -33 110
rect 33 84 63 110
rect 129 84 159 110
rect -159 -110 -129 -84
rect -63 -110 -33 -84
rect 33 -110 63 -84
rect 129 -110 159 -84
<< locali >>
rect -323 233 -227 267
rect 227 233 323 267
rect -323 171 -289 233
rect 289 171 323 233
rect -209 72 -175 88
rect -209 -88 -175 -72
rect -113 72 -79 88
rect -113 -88 -79 -72
rect -17 72 17 88
rect -17 -88 17 -72
rect 79 72 113 88
rect 79 -88 113 -72
rect 175 72 209 88
rect 175 -88 209 -72
rect -323 -233 -289 -171
rect 289 -233 323 -171
<< viali >>
rect -209 -72 -175 72
rect -113 -72 -79 72
rect -17 -72 17 72
rect 79 -72 113 72
rect 175 -72 209 72
<< metal1 >>
rect -215 72 -169 84
rect -215 -72 -209 72
rect -175 -72 -169 72
rect -215 -84 -169 -72
rect -119 72 -73 84
rect -119 -72 -113 72
rect -79 -72 -73 72
rect -119 -84 -73 -72
rect -23 72 23 84
rect -23 -72 -17 72
rect 17 -72 23 72
rect -23 -84 23 -72
rect 73 72 119 84
rect 73 -72 79 72
rect 113 -72 119 72
rect 73 -84 119 -72
rect 169 72 215 84
rect 169 -72 175 72
rect 209 -72 215 72
rect 169 -84 215 -72
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -306 -250 306 250
string parameters w 0.84 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
