**.subckt tb_charge_pump
VSS vss GND {vss} 
VDD vdd vss {vdd} 
Vref net2 vss PULSE(0 {vin} 0 1p 1p {Tref/2} {Tref}) DC {vin} AC 0 
Vdiv net1 vss PULSE(0 {vin} 0 1p 1p {Tref/2} {Tref}) DC {vin} AC 0 
C1 net3 vss 33.5p m=1
R1 vctrl net3 2k m=1
C2 vctrl vss 6.7p m=1
vout cp_out vctrl 0
x1 vss vdd net16 net17 net18 net19 Reset PFD
x5 vdd net4 net2 vss inverter_cp_x2
x6 vdd QA net4 vss inverter_cp_x2
x7 vdd net5 net1 vss inverter_cp_x2
x8 vdd QB net5 vss inverter_cp_x2
x3 Up vdd QA nUp Down QB vss nDown pfd_cp_interface_pex_c
x2 vdd Up nUp cp_out Down nDown vss iref_cp nswitch pswitch biasp charge_pump_pex_c
I0 net6 vss 100u
x4 vdd net6 vss iref_cp net7 net8 net9 net10 net11 net12 net13 net14 net15 bias_pex_c
**** begin user architecture code



* Parameters
.param kp = 1.0
.param vdd = kp*1.8
.param vss = 0.0
.param vin = vdd
.param fref = 100e6
.param Tref = 1/fref
.param Cn = 0.0001fF
.param Cp = 0.0001fF
.param iref=100u

.options TEMP = 100.0
.options RSHUNT = 1e20

* Models
.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib SS
*.include ~/caravel_analog_fulgor/xschem/simulations/simulations/PFD_pex_c.spice
.include ~/caravel_analog_fulgor/xschem/simulations/pfd_cp_interface_pex_c.spice
.include ~/caravel_analog_fulgor/xschem/simulations/charge_pump_pex_c.spice
.include ~/caravel_analog_fulgor/xschem/simulations/bias_pex_c.spice

* Data to save
.save all

.ic v(A) = 0.0
.ic v(B) = 0.0
.ic v(vctrl) = 0.0

* Simulation
.control
	op
	echo .
	echo ---- M1 bias ----
	print @M.X4.XM1.msky130_fd_pr__pfet_01v8_lvt[id]
	print @M.X4.XM1.msky130_fd_pr__pfet_01v8_lvt[vds]
	print @M.X4.XM1.msky130_fd_pr__pfet_01v8_lvt[vdsat]
	print @M.X4.XM1.msky130_fd_pr__pfet_01v8_lvt[vgs]
	echo ---- M2 bias ----
	print @M.X4.XM2.msky130_fd_pr__pfet_01v8_lvt[id]
	print @M.X4.XM2.msky130_fd_pr__pfet_01v8_lvt[vds]
	print @M.X4.XM2.msky130_fd_pr__pfet_01v8_lvt[vdsat]
	print @M.X4.XM2.msky130_fd_pr__pfet_01v8_lvt[vgs]
	echo ---- M3 bias ----
	print @M.X4.XM3.msky130_fd_pr__pfet_01v8_lvt[id]
	print @M.X4.XM3.msky130_fd_pr__pfet_01v8_lvt[vds]
	print @M.X4.XM3.msky130_fd_pr__pfet_01v8_lvt[vdsat]
	print @M.X4.XM3.msky130_fd_pr__pfet_01v8_lvt[vgs]
	echo ---- M4 bias ----
	print @M.X4.XM4.msky130_fd_pr__pfet_01v8_lvt[id]
	print @M.X4.XM4.msky130_fd_pr__pfet_01v8_lvt[vds]
	print @M.X4.XM4.msky130_fd_pr__pfet_01v8_lvt[vdsat]
	print @M.X4.XM4.msky130_fd_pr__pfet_01v8_lvt[vgs]
	echo ---- M5 bias ----
	print @M.X4.XM5.msky130_fd_pr__nfet_01v8[id]
	print @M.X4.XM5.msky130_fd_pr__nfet_01v8[vds]
	print @M.X4.XM5.msky130_fd_pr__nfet_01v8[vdsat]
	print @M.X4.XM5.msky130_fd_pr__nfet_01v8[vgs]
	echo ---- M6 bias ----
	print @M.X4.XM6.msky130_fd_pr__nfet_01v8[id]
	print @M.X4.XM6.msky130_fd_pr__nfet_01v8[vds]
	print @M.X4.XM6.msky130_fd_pr__nfet_01v8[vdsat]
	print @M.X4.XM6.msky130_fd_pr__nfet_01v8[vgs]
	echo ---- M7 bias ----
	print @M.X4.XM7.msky130_fd_pr__pfet_01v8[id]
	print @M.X4.XM7.msky130_fd_pr__pfet_01v8[vds]
	print @M.X4.XM7.msky130_fd_pr__pfet_01v8[vdsat]
	print @M.X4.XM7.msky130_fd_pr__pfet_01v8[vgs]
	echo --- Cgs ---
	print @M.X2.XM7.msky130_fd_pr__pfet_01v8[cgs]
	print @M.X2.XM8.msky130_fd_pr__nfet_01v8[cgs]
	echo --- Cgs ---
	print @M.X2.XM7.msky130_fd_pr__pfet_01v8[cgd]
	print @M.X2.XM8.msky130_fd_pr__nfet_01v8[cgd]
	echo --- Cgs ---
	print @M.X2.XM7.msky130_fd_pr__pfet_01v8[cgb]
	print @M.X2.XM8.msky130_fd_pr__nfet_01v8[cgb]
	echo --- Cgs ---
	print @M.X2.XM7.msky130_fd_pr__pfet_01v8[cgg]
	print @M.X2.XM8.msky130_fd_pr__nfet_01v8[cgg]

	reset


	tran 0.01ns 400ns
	write tb_cp_gate_switched_tran.raw
	plot i(v.x2.vm1) i(v.x2.vm2)
	plot v(vctrl) v(nDown)+2 v(Down)+4 v(nUp)+6 v(Up)+8 v(QB)+10 v(QA)+12
	plot v(pswitch) v(nswitch) xlimit 4ns 44ns
.endc



**** end user architecture code
**.ends

* expanding   symbol:  PFD.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/PFD.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/PFD.sch
.subckt PFD  vss vdd Up A B Down Reset
*.iopin vdd
*.iopin vss
*.ipin A
*.ipin B
*.opin Down
*.opin Up
*.iopin Reset
x1 vdd A Up Reset vss DFF
x2 vdd B Down Reset vss DFF
x3 vdd Reset Up Down vss and_pfd
.ends


* expanding   symbol:  inverter_cp_x2.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_cp_x2.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_cp_x2.sch
.subckt inverter_cp_x2  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
.ends


* expanding   symbol:  DFF.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/DFF.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/DFF.sch
.subckt DFF  D CLK Q Reset vss
*.ipin D
*.ipin CLK
*.opin Q
*.ipin Reset
*.iopin vss
x1 D CLK Q P vss nor
x2 D P P1 Q vss nor
x3 D P P2 P1 vss nor
x4 D P1 Reset P2 vss nor
.ends


* expanding   symbol:  and_pfd.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/and_pfd.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/and_pfd.sch
.subckt and_pfd  vdd out A B vss
*.iopin vdd
*.iopin vss
*.opin out
*.ipin A
*.ipin B
XM1 out_nand A net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out_nand A vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net1 B vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 out_nand B net2 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 net2 A vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 out_nand B vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 out out_nand vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 out out_nand vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  nor.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/nor.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/nor.sch
.subckt nor  vdd A B out vss
*.ipin A
*.ipin B
*.iopin vdd
*.opin out
*.iopin vss
XM1 out A vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out B vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 out B net1 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net1 A vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 net2 B vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 out A net2 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

.GLOBAL GND
** flattened .save nodes
.end
