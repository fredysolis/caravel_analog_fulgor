**.subckt cap3_loop_filter in out
*.iopin in
*.iopin out
XC1 in out sky130_fd_pr__cap_mim_m3_1 W=20 L=20 MF=4 m=4
**.ends
** flattened .save nodes
.end
