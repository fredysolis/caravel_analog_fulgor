magic
tech sky130A
magscale 1 2
timestamp 1624896651
<< nwell >>
rect 2984 3068 4571 3079
rect 10778 3059 11706 3083
<< metal1 >>
rect -1746 6066 36 6106
rect -1746 6012 149 6066
rect -1746 5972 36 6012
rect -1745 3883 -1188 5972
rect 17525 5699 17853 5700
rect 17525 5692 21244 5699
rect 17525 5376 20937 5692
rect 21232 5376 21244 5692
rect 17525 5371 21244 5376
rect 11727 5280 11848 5293
rect 11676 5120 11686 5280
rect 11841 5120 11851 5280
rect 11727 5098 11848 5120
rect 17525 4766 17853 5371
rect 19149 5370 21244 5371
rect 18332 4902 18342 4981
rect 18516 4902 18526 4981
rect 18760 4902 19117 4982
rect 19474 4903 19484 4988
rect 19645 4903 19655 4988
rect 11366 4438 17853 4766
rect 14091 3992 16674 4150
rect 1 3108 11416 3119
rect 1 3099 11506 3108
rect 0 3037 11506 3099
rect 1 3031 11506 3037
rect 1 3013 11416 3031
rect 2870 2904 11416 3013
rect 14091 2792 14249 3992
rect 16516 2950 16674 3992
rect 18812 2983 19229 4339
rect 21313 4070 23316 4148
rect 21313 3992 22312 4070
rect 21313 2923 21471 3992
rect -1702 1698 -1395 2597
rect 14346 2347 14356 2506
rect 14531 2347 14541 2506
rect 15177 1698 15539 2757
rect 21597 2241 21607 2338
rect 21754 2241 21764 2338
rect -1702 1370 391 1698
rect 14120 1370 16525 1698
rect 20954 1438 20964 1663
rect 21241 1438 21251 1663
rect -1702 1181 -1395 1370
rect 22532 1369 22819 2760
rect 21748 1270 22932 1369
rect 21748 1204 22896 1270
rect 22532 1196 22819 1204
rect -1948 673 -1938 743
rect -1688 673 -1678 743
rect -1425 674 -1415 741
rect -1213 674 -1203 741
rect 22373 672 22383 740
rect 22535 672 22545 740
rect 22817 678 22827 740
rect 22968 678 22978 740
rect -1329 94 86 134
rect -1351 40 101 94
rect -1326 30 86 40
rect 14232 30 16473 164
rect 21723 143 22442 179
rect 21742 138 22442 143
rect 21707 84 22470 138
rect 21745 80 22442 84
rect 21679 44 22442 80
<< via1 >>
rect 20937 5376 21232 5692
rect 11686 5120 11841 5280
rect 18342 4902 18516 4981
rect 19484 4903 19645 4988
rect 14356 2347 14531 2506
rect 21607 2241 21754 2338
rect 20964 1438 21241 1663
rect -1938 673 -1688 743
rect -1415 674 -1213 741
rect 22383 672 22535 740
rect 22827 678 22968 740
<< metal2 >>
rect 20937 5692 21232 5702
rect 20937 5366 21232 5376
rect 11686 5280 11841 5290
rect 15870 5265 15968 5272
rect 11841 5262 15970 5265
rect 11841 5138 15870 5262
rect 15968 5138 15970 5262
rect 11841 5135 15970 5138
rect 15870 5128 15968 5135
rect 11686 5110 11841 5120
rect 23186 5013 23271 5016
rect 19564 5007 23271 5013
rect 19564 4998 23186 5007
rect 16085 4989 16196 4998
rect 19484 4991 23186 4998
rect 18342 4989 18516 4991
rect 16082 4988 18522 4989
rect 16082 4897 16085 4988
rect 16196 4981 18522 4988
rect 16196 4902 18342 4981
rect 18516 4902 18522 4981
rect 16196 4897 18522 4902
rect 19479 4988 23186 4991
rect 19479 4903 19484 4988
rect 19645 4903 23186 4988
rect 19479 4899 23186 4903
rect 18342 4892 18516 4897
rect 19484 4895 23186 4899
rect 23271 4899 23273 4991
rect 19484 4893 23271 4895
rect 16085 4876 16196 4886
rect 19564 4885 23271 4893
rect 22884 3484 22975 3494
rect 15070 3470 15167 3480
rect 15070 3367 15167 3377
rect 15570 3473 15667 3483
rect 15570 3370 15667 3380
rect 22384 3473 22468 3483
rect 22384 3374 22468 3384
rect 22884 3373 22975 3383
rect -1394 3237 -1242 3247
rect -1951 3151 -1763 3161
rect -1394 3118 -1242 3128
rect 16084 3101 16193 3108
rect -1951 3061 -1763 3071
rect 15338 3098 16196 3101
rect -2235 2687 -2151 2980
rect -972 2687 -876 2980
rect 15338 2857 16084 3098
rect 16193 2857 16196 3098
rect 15338 2856 16196 2857
rect 16084 2847 16193 2856
rect 22635 2841 22727 3134
rect 14356 2506 14531 2516
rect 14765 2506 14864 2514
rect 14531 2504 14864 2506
rect 14531 2351 14765 2504
rect 14531 2347 14864 2351
rect 22085 2348 22166 2356
rect 14356 2337 14531 2347
rect 14765 2341 14864 2347
rect 21599 2346 22170 2348
rect 21599 2338 22085 2346
rect 21599 2241 21607 2338
rect 21754 2241 22085 2338
rect 21599 2235 22085 2241
rect 22166 2235 22170 2346
rect 21599 2231 22170 2235
rect 22085 2225 22166 2231
rect 20964 1663 21241 1673
rect 20964 1428 21241 1438
rect -1938 743 -1688 753
rect -1938 663 -1688 673
rect -1415 741 -1213 751
rect -1415 664 -1213 674
rect 22383 740 22535 750
rect 22383 662 22535 672
rect 22827 740 22968 750
rect 22827 668 22968 678
<< via2 >>
rect 20937 5376 21232 5692
rect 15870 5138 15968 5262
rect 16085 4886 16196 4988
rect 23186 4895 23271 5007
rect 15070 3377 15167 3470
rect 15570 3380 15667 3473
rect 22384 3384 22468 3473
rect 22884 3383 22975 3484
rect -1951 3071 -1763 3151
rect -1394 3128 -1242 3237
rect 16084 2857 16193 3098
rect 14765 2351 14864 2504
rect 22085 2235 22166 2346
rect 20964 1438 21241 1663
rect -1938 673 -1688 743
rect -1415 674 -1213 741
rect 22383 672 22535 740
rect 22827 678 22968 740
<< metal3 >>
rect 20927 5692 21242 5697
rect 20927 5376 20937 5692
rect 21232 5376 21242 5692
rect 20927 5371 21242 5376
rect -2788 5275 -2700 5279
rect -2792 5185 -2786 5275
rect -2701 5185 -2691 5275
rect 15860 5262 15978 5267
rect -2788 3566 -2700 5185
rect 15860 5138 15870 5262
rect 15968 5138 15978 5262
rect 15860 5133 15978 5138
rect -1518 4023 -1430 4026
rect -1527 3933 -1517 4023
rect -1431 3933 -1421 4023
rect -1676 3623 -1608 3769
rect -2780 3485 -2710 3566
rect -1961 3151 -1753 3156
rect -1961 3071 -1951 3151
rect -1763 3071 -1753 3151
rect -1961 3066 -1753 3071
rect -1941 748 -1853 3066
rect -1686 953 -1598 3623
rect -1518 3594 -1430 3933
rect 14780 3791 14850 3934
rect -402 3696 -334 3769
rect -1510 3486 -1440 3594
rect -1404 3237 -1210 3242
rect -1404 3128 -1394 3237
rect -1242 3128 -1210 3237
rect -1404 3123 -1210 3128
rect -1695 879 -1685 953
rect -1599 879 -1589 953
rect -1686 875 -1598 879
rect -1948 743 -1678 748
rect -1298 746 -1210 3123
rect -412 2189 -324 3696
rect 14772 2509 14860 3791
rect 15874 3739 15962 5133
rect 16075 4988 16206 4993
rect 16075 4886 16085 4988
rect 16196 4886 16206 4988
rect 16075 4881 16206 4886
rect 15884 3640 15954 3739
rect 15074 3475 15162 3493
rect 15572 3478 15660 3481
rect 15060 3470 15177 3475
rect 15060 3377 15070 3470
rect 15167 3377 15177 3470
rect 15060 3372 15177 3377
rect 15560 3473 15677 3478
rect 15560 3380 15570 3473
rect 15667 3380 15677 3473
rect 15560 3375 15677 3380
rect 14755 2504 14874 2509
rect 14755 2351 14765 2504
rect 14864 2351 14874 2504
rect 14755 2346 14874 2351
rect -421 2115 -411 2189
rect -325 2115 -315 2189
rect -412 2114 -324 2115
rect -1948 673 -1938 743
rect -1688 673 -1678 743
rect -1948 668 -1678 673
rect -1425 741 -1203 746
rect -1425 674 -1415 741
rect -1213 674 -1203 741
rect -1425 669 -1203 674
rect -1941 373 -1853 668
rect -1307 630 -1203 669
rect 15074 631 15162 3372
rect -1307 511 -1297 630
rect -1210 511 -1200 630
rect -1298 509 -1210 511
rect 15064 508 15074 631
rect 15162 508 15172 631
rect 15074 501 15162 508
rect -1962 237 -1952 373
rect -1845 237 -1835 373
rect 15572 363 15660 3375
rect 16081 3103 16198 4881
rect 16074 3098 16203 3103
rect 16074 2857 16084 3098
rect 16193 2857 16203 3098
rect 16074 2852 16203 2857
rect 16081 1609 16198 2852
rect 20986 1668 21183 5371
rect 23184 5012 23272 5016
rect 23176 5007 23281 5012
rect 23176 4895 23186 5007
rect 23271 4895 23281 5007
rect 23176 4890 23281 4895
rect 22090 3817 22160 3967
rect 22082 2351 22170 3817
rect 23184 3749 23272 4890
rect 23194 3640 23264 3749
rect 22381 3478 22469 3487
rect 22874 3484 22985 3489
rect 22374 3473 22478 3478
rect 22374 3384 22384 3473
rect 22468 3384 22478 3473
rect 22374 3379 22478 3384
rect 22874 3383 22884 3484
rect 22975 3383 22985 3484
rect 22075 2346 22176 2351
rect 22075 2235 22085 2346
rect 22166 2235 22176 2346
rect 22075 2230 22176 2235
rect 22082 2224 22170 2230
rect 20954 1663 21251 1668
rect 16081 1492 16598 1609
rect 20954 1438 20964 1663
rect 21241 1438 21251 1663
rect 20954 1433 21251 1438
rect 22381 745 22469 3379
rect 22874 3378 22985 3383
rect 22882 745 22970 3378
rect 22373 740 22545 745
rect 22373 672 22383 740
rect 22535 672 22545 740
rect 22817 740 22978 745
rect 22817 678 22827 740
rect 22968 678 22978 740
rect 22817 673 22978 678
rect 22373 667 22545 672
rect 15562 240 15572 363
rect 15660 240 15670 363
<< via3 >>
rect -2786 5185 -2701 5275
rect -1517 3933 -1431 4023
rect -1685 879 -1599 953
rect -411 2115 -325 2189
rect -1297 511 -1210 630
rect 15074 508 15162 631
rect -1952 237 -1845 373
rect 15572 240 15660 363
<< metal4 >>
rect -2792 5275 2396 5276
rect -2792 5185 -2786 5275
rect -2701 5185 2396 5275
rect -2792 5184 2396 5185
rect -1522 4023 2450 4024
rect -1522 3933 -1517 4023
rect -1431 3933 2450 4023
rect -1522 3932 2450 3933
rect -412 2189 -324 2190
rect -412 2115 -411 2189
rect -325 2185 -324 2189
rect -325 2119 2959 2185
rect -325 2115 -324 2119
rect -412 2114 -324 2115
rect -1686 953 -1598 954
rect -1686 879 -1685 953
rect -1599 949 -1598 953
rect -1599 883 2950 949
rect -1599 879 -1598 883
rect -1686 878 -1598 879
rect 15073 631 15163 632
rect -1298 630 15074 631
rect -1298 511 -1297 630
rect -1210 511 15074 630
rect -1298 510 15074 511
rect -1296 508 15074 510
rect 15162 508 15172 631
rect 15073 507 15163 508
rect -1953 373 -1844 374
rect -1953 237 -1952 373
rect -1845 363 -1844 373
rect 15571 363 15661 364
rect -1845 240 15572 363
rect 15660 240 15661 363
rect -1845 237 -1844 240
rect 15571 239 15661 240
rect -1953 236 -1844 237
use div_by_5  div_by_5_0
timestamp 1624896651
transform 1 0 556 0 1 0
box -556 0 13892 3068
use div_by_2  div_by_2_0
timestamp 1624896651
transform 1 0 17530 0 1 0
box -1244 0 4228 3068
use mux2to1  mux2to1_1
timestamp 1624653480
transform -1 0 23305 0 -1 2710
box -11 -1360 1267 2
use mux2to1  mux2to1_0
timestamp 1624653480
transform -1 0 15995 0 -1 2710
box -11 -1360 1267 2
use mux2to4  mux2to4_0
timestamp 1624653480
transform 1 0 -2821 0 -1 2556
box -11 -1360 2541 2
use inverter_min_x2  inverter_min_x2_2
timestamp 1624049879
transform 1 0 -1766 0 -1 655
box -53 -615 473 655
use inverter_min_x2  inverter_min_x2_1
timestamp 1624049879
transform -1 0 22879 0 -1 655
box -53 -615 473 655
use inverter_min_x4  inverter_min_x4_0
timestamp 1624049879
transform 1 0 18971 0 -1 4889
box -53 -616 665 643
use inverter_min_x2  inverter_min_x2_0
timestamp 1624049879
transform 1 0 18445 0 -1 4890
box -53 -615 473 655
use prescaler_23  prescaler_23_0
timestamp 1624896651
transform 1 0 0 0 -1 6136
box 0 -316 11752 3068
<< labels >>
rlabel metal2 22635 2841 22727 3134 1 out
rlabel metal4 -2701 5184 2396 5276 1 clk_0
rlabel metal4 -1431 3932 2450 4024 1 n_clk_0
rlabel metal4 -325 2119 2959 2185 1 n_clk_1
rlabel metal4 -1599 883 2950 949 1 clk_1
rlabel metal2 14531 2347 14765 2506 1 clk_5
rlabel metal2 11841 5135 15870 5265 1 clk_pre
rlabel metal2 19645 4885 23186 5013 1 clk_d
rlabel metal2 21754 2231 22085 2348 1 clk_2
rlabel metal3 16081 3098 16198 4886 1 clk_out_mux21
rlabel metal3 22882 740 22970 3383 1 s_1
rlabel metal3 22381 740 22469 3384 1 s_1_n
rlabel metal3 -1941 373 -1853 673 1 s_0
rlabel metal3 -1307 630 -1203 674 1 s_0_n
rlabel metal1 14232 30 16473 164 1 vdd
rlabel metal1 19149 5370 20937 5699 1 vss
rlabel metal2 -972 2687 -876 2980 1 in_b
rlabel metal2 -2235 2687 -2151 2980 1 in_a
<< end >>
