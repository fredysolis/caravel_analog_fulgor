* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_4798MH VSUBS a_81_n156# a_111_n125# a_15_n125# a_n173_n125#
+ w_n311_n344# a_n111_n156# a_n15_n156# a_n81_n125#
X0 a_n81_n125# a_n111_n156# a_n173_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n15_n156# a_n81_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_81_n156# a_15_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n81_n125# w_n311_n344# 0.09fF
C1 a_n15_n156# a_81_n156# 0.02fF
C2 w_n311_n344# a_n173_n125# 0.14fF
C3 a_15_n125# w_n311_n344# 0.09fF
C4 a_n81_n125# a_n173_n125# 0.36fF
C5 a_111_n125# w_n311_n344# 0.14fF
C6 a_n81_n125# a_15_n125# 0.36fF
C7 a_n81_n125# a_111_n125# 0.13fF
C8 a_n111_n156# a_n15_n156# 0.02fF
C9 a_15_n125# a_n173_n125# 0.13fF
C10 a_111_n125# a_n173_n125# 0.08fF
C11 a_15_n125# a_111_n125# 0.36fF
C12 a_111_n125# VSUBS 0.03fF
C13 a_15_n125# VSUBS 0.03fF
C14 a_n81_n125# VSUBS 0.03fF
C15 a_n173_n125# VSUBS 0.03fF
C16 a_81_n156# VSUBS 0.05fF
C17 a_n15_n156# VSUBS 0.05fF
C18 a_n111_n156# VSUBS 0.05fF
C19 w_n311_n344# VSUBS 2.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_BHR94T a_n15_n151# w_n311_n335# a_81_n151# a_111_n125#
+ a_15_n125# a_n173_n125# a_n111_n151# a_n81_n125#
X0 a_111_n125# a_81_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n15_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n111_n151# a_n15_n151# 0.02fF
C1 a_n173_n125# a_111_n125# 0.08fF
C2 a_n15_n151# a_81_n151# 0.02fF
C3 a_n173_n125# a_n81_n125# 0.36fF
C4 a_n81_n125# a_111_n125# 0.13fF
C5 a_n173_n125# a_15_n125# 0.13fF
C6 a_15_n125# a_111_n125# 0.36fF
C7 a_n81_n125# a_15_n125# 0.36fF
C8 a_111_n125# w_n311_n335# 0.17fF
C9 a_15_n125# w_n311_n335# 0.12fF
C10 a_n81_n125# w_n311_n335# 0.12fF
C11 a_n173_n125# w_n311_n335# 0.17fF
C12 a_81_n151# w_n311_n335# 0.05fF
C13 a_n15_n151# w_n311_n335# 0.05fF
C14 a_n111_n151# w_n311_n335# 0.05fF
.ends

.subckt trans_gate m1_187_n605# vss m1_45_n513# vdd
Xsky130_fd_pr__pfet_01v8_4798MH_0 vss vss m1_187_n605# m1_45_n513# m1_45_n513# vdd
+ vss vss m1_187_n605# sky130_fd_pr__pfet_01v8_4798MH
Xsky130_fd_pr__nfet_01v8_BHR94T_0 vdd vss vdd m1_187_n605# m1_45_n513# m1_45_n513#
+ vdd m1_187_n605# sky130_fd_pr__nfet_01v8_BHR94T
C0 m1_187_n605# vdd 0.55fF
C1 m1_45_n513# vdd 0.69fF
C2 m1_45_n513# m1_187_n605# 0.36fF
C3 m1_187_n605# vss 0.93fF
C4 m1_45_n513# vss 1.31fF
C5 vdd vss 3.36fF
.ends

.subckt sky130_fd_pr__pfet_01v8_7KT7MH VSUBS a_n111_n186# a_111_n125# a_15_n125# a_n173_n125#
+ w_n311_n344# a_n81_n125#
X0 a_n81_n125# a_n111_n186# a_n173_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n111_n186# a_n81_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_n111_n186# a_15_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_15_n125# a_n173_n125# 0.13fF
C1 w_n311_n344# a_n81_n125# 0.09fF
C2 a_15_n125# w_n311_n344# 0.09fF
C3 w_n311_n344# a_n173_n125# 0.14fF
C4 a_n81_n125# a_111_n125# 0.13fF
C5 a_15_n125# a_111_n125# 0.36fF
C6 a_n173_n125# a_111_n125# 0.08fF
C7 w_n311_n344# a_111_n125# 0.14fF
C8 a_15_n125# a_n81_n125# 0.36fF
C9 a_n81_n125# a_n173_n125# 0.36fF
C10 a_111_n125# VSUBS 0.03fF
C11 a_15_n125# VSUBS 0.03fF
C12 a_n81_n125# VSUBS 0.03fF
C13 a_n173_n125# VSUBS 0.03fF
C14 a_n111_n186# VSUBS 0.26fF
C15 w_n311_n344# VSUBS 2.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS6QM w_n311_n335# a_111_n125# a_15_n125# a_n173_n125#
+ a_n111_n151# a_n81_n125#
X0 a_111_n125# a_n111_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n111_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_111_n125# a_n81_n125# 0.13fF
C1 a_15_n125# a_n173_n125# 0.13fF
C2 a_111_n125# a_n173_n125# 0.08fF
C3 a_n81_n125# a_n173_n125# 0.36fF
C4 a_111_n125# a_15_n125# 0.36fF
C5 a_15_n125# a_n81_n125# 0.36fF
C6 a_111_n125# w_n311_n335# 0.17fF
C7 a_15_n125# w_n311_n335# 0.12fF
C8 a_n81_n125# w_n311_n335# 0.12fF
C9 a_n173_n125# w_n311_n335# 0.17fF
C10 a_n111_n151# w_n311_n335# 0.25fF
.ends

.subckt inverter_cp_x1 out in vss vdd
Xsky130_fd_pr__pfet_01v8_7KT7MH_0 vss in out vdd vdd vdd out sky130_fd_pr__pfet_01v8_7KT7MH
Xsky130_fd_pr__nfet_01v8_2BS6QM_0 vss out vss vss in out sky130_fd_pr__nfet_01v8_2BS6QM
C0 out in 0.32fF
C1 out vdd 0.10fF
C2 out vss 0.77fF
C3 in vss 0.95fF
C4 vdd vss 3.13fF
.ends

.subckt clock_inverter vss inverter_cp_x1_2/in CLK vdd inverter_cp_x1_0/out CLK_d
+ nCLK_d
Xtrans_gate_0 nCLK_d vss inverter_cp_x1_0/out vdd trans_gate
Xinverter_cp_x1_0 inverter_cp_x1_0/out CLK vss vdd inverter_cp_x1
Xinverter_cp_x1_2 CLK_d inverter_cp_x1_2/in vss vdd inverter_cp_x1
Xinverter_cp_x1_1 inverter_cp_x1_2/in CLK vss vdd inverter_cp_x1
C0 vdd inverter_cp_x1_2/in 0.21fF
C1 CLK inverter_cp_x1_2/in 0.31fF
C2 inverter_cp_x1_0/out vdd 0.28fF
C3 CLK_d inverter_cp_x1_2/in 0.12fF
C4 vdd CLK 0.36fF
C5 nCLK_d vdd 0.03fF
C6 inverter_cp_x1_0/out CLK 0.31fF
C7 CLK_d vdd 0.03fF
C8 nCLK_d inverter_cp_x1_0/out 0.11fF
C9 inverter_cp_x1_2/in vss 2.01fF
C10 CLK_d vss 0.96fF
C11 inverter_cp_x1_0/out vss 1.97fF
C12 CLK vss 3.03fF
C13 vdd vss 16.51fF
C14 nCLK_d vss 1.44fF
.ends

.subckt sky130_fd_pr__pfet_01v8_MJG8BZ VSUBS a_n125_n95# a_63_n95# w_n263_n314# a_n33_n95#
+ a_n63_n192#
X0 a_63_n95# a_n63_n192# a_n33_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n33_n95# a_n63_n192# a_n125_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
C0 a_n125_n95# w_n263_n314# 0.11fF
C1 a_n125_n95# a_63_n95# 0.10fF
C2 a_n125_n95# a_n33_n95# 0.28fF
C3 w_n263_n314# a_63_n95# 0.11fF
C4 w_n263_n314# a_n33_n95# 0.08fF
C5 a_63_n95# a_n33_n95# 0.28fF
C6 a_63_n95# VSUBS 0.03fF
C7 a_n33_n95# VSUBS 0.03fF
C8 a_n125_n95# VSUBS 0.03fF
C9 a_n63_n192# VSUBS 0.20fF
C10 w_n263_n314# VSUBS 1.80fF
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS854 w_n311_n335# a_n129_n213# a_111_n125# a_15_n125#
+ a_n173_n125# a_n81_n125#
X0 a_111_n125# a_n129_n213# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n129_n213# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n129_n213# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n81_n125# a_n173_n125# 0.36fF
C1 a_n173_n125# a_n129_n213# 0.02fF
C2 a_n173_n125# a_111_n125# 0.08fF
C3 a_n173_n125# a_15_n125# 0.13fF
C4 a_n81_n125# a_n129_n213# 0.10fF
C5 a_n81_n125# a_111_n125# 0.13fF
C6 a_n81_n125# a_15_n125# 0.36fF
C7 a_n129_n213# a_111_n125# 0.01fF
C8 a_n129_n213# a_15_n125# 0.10fF
C9 a_111_n125# a_15_n125# 0.36fF
C10 a_111_n125# w_n311_n335# 0.05fF
C11 a_15_n125# w_n311_n335# 0.05fF
C12 a_n81_n125# w_n311_n335# 0.05fF
C13 a_n173_n125# w_n311_n335# 0.05fF
C14 a_n129_n213# w_n311_n335# 0.49fF
.ends

.subckt sky130_fd_pr__nfet_01v8_KU9PSX a_n125_n95# a_n33_n95# a_n81_n183# w_n263_n305#
X0 a_n33_n95# a_n81_n183# a_n125_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n125_n95# a_n81_n183# a_n33_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
C0 a_n33_n95# a_n125_n95# 0.88fF
C1 a_n125_n95# a_n81_n183# 0.16fF
C2 a_n33_n95# a_n81_n183# 0.10fF
C3 a_n33_n95# w_n263_n305# 0.07fF
C4 a_n125_n95# w_n263_n305# 0.13fF
C5 a_n81_n183# w_n263_n305# 0.31fF
.ends

.subckt latch_diff m1_657_280# nQ Q vss CLK vdd nD D
Xsky130_fd_pr__pfet_01v8_MJG8BZ_0 vss vdd vdd vdd nQ Q sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__pfet_01v8_MJG8BZ_1 vss vdd vdd vdd Q nQ sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__nfet_01v8_2BS854_0 vss CLK vss m1_657_280# m1_657_280# vss sky130_fd_pr__nfet_01v8_2BS854
Xsky130_fd_pr__nfet_01v8_KU9PSX_0 m1_657_280# Q nD vss sky130_fd_pr__nfet_01v8_KU9PSX
Xsky130_fd_pr__nfet_01v8_KU9PSX_1 m1_657_280# nQ D vss sky130_fd_pr__nfet_01v8_KU9PSX
C0 nQ D 0.05fF
C1 m1_657_280# nQ 1.41fF
C2 vdd nQ 0.16fF
C3 nD Q 0.05fF
C4 Q D 0.05fF
C5 m1_657_280# Q 0.94fF
C6 vdd Q 0.16fF
C7 nQ Q 0.93fF
C8 nD nQ 0.05fF
C9 m1_657_280# CLK 0.24fF
C10 D vss 0.53fF
C11 Q vss -0.55fF
C12 m1_657_280# vss 1.88fF
C13 nD vss 0.16fF
C14 CLK vss 0.87fF
C15 nQ vss 1.16fF
C16 vdd vss 5.98fF
.ends

.subckt DFlipFlop latch_diff_0/m1_657_280# vss vdd latch_diff_1/D clock_inverter_0/inverter_cp_x1_2/in
+ nQ nCLK latch_diff_0/nD Q latch_diff_1/nD latch_diff_1/m1_657_280# D latch_diff_0/D
+ CLK clock_inverter_0/inverter_cp_x1_0/out
Xclock_inverter_0 vss clock_inverter_0/inverter_cp_x1_2/in D vdd clock_inverter_0/inverter_cp_x1_0/out
+ latch_diff_0/D latch_diff_0/nD clock_inverter
Xlatch_diff_0 latch_diff_0/m1_657_280# latch_diff_1/nD latch_diff_1/D vss CLK vdd
+ latch_diff_0/nD latch_diff_0/D latch_diff
Xlatch_diff_1 latch_diff_1/m1_657_280# nQ Q vss nCLK vdd latch_diff_1/nD latch_diff_1/D
+ latch_diff
C0 vdd clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C1 latch_diff_1/D latch_diff_0/m1_657_280# 0.43fF
C2 latch_diff_0/nD vdd 0.14fF
C3 latch_diff_1/m1_657_280# latch_diff_1/nD 0.42fF
C4 latch_diff_0/nD latch_diff_1/D 0.41fF
C5 nQ latch_diff_1/nD 0.08fF
C6 latch_diff_0/nD latch_diff_0/m1_657_280# 0.38fF
C7 latch_diff_1/m1_657_280# latch_diff_1/D 0.32fF
C8 latch_diff_0/D latch_diff_1/nD 0.04fF
C9 latch_diff_1/D nQ 0.11fF
C10 latch_diff_1/m1_657_280# latch_diff_0/m1_657_280# 0.18fF
C11 Q latch_diff_1/nD 0.01fF
C12 vdd latch_diff_0/D 0.09fF
C13 latch_diff_1/D latch_diff_0/D 0.11fF
C14 vdd latch_diff_1/nD 0.02fF
C15 latch_diff_0/m1_657_280# latch_diff_0/D 0.37fF
C16 latch_diff_1/D latch_diff_1/nD 0.33fF
C17 latch_diff_0/m1_657_280# latch_diff_1/nD 0.14fF
C18 vdd latch_diff_1/D 0.03fF
C19 Q vss -0.92fF
C20 latch_diff_1/m1_657_280# vss 0.64fF
C21 nCLK vss 0.83fF
C22 nQ vss 0.57fF
C23 latch_diff_1/D vss -0.30fF
C24 latch_diff_0/m1_657_280# vss 0.72fF
C25 CLK vss 0.83fF
C26 latch_diff_1/nD vss 1.83fF
C27 clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C28 latch_diff_0/D vss 1.29fF
C29 clock_inverter_0/inverter_cp_x1_0/out vss 1.84fF
C30 D vss 3.27fF
C31 vdd vss 32.62fF
C32 latch_diff_0/nD vss 1.74fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ZP3U9B VSUBS a_n221_n84# a_159_n84# w_n359_n303# a_n63_n110#
+ a_n129_n84# a_33_n110# a_n159_n110# a_63_n84# a_129_n110# a_n33_n84#
X0 a_n129_n84# a_n159_n110# a_n221_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_63_n84# a_33_n110# a_n33_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_n33_n84# a_n63_n110# a_n129_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_159_n84# a_129_n110# a_63_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 w_n359_n303# a_n129_n84# 0.06fF
C1 w_n359_n303# a_159_n84# 0.08fF
C2 w_n359_n303# a_n221_n84# 0.08fF
C3 w_n359_n303# a_n33_n84# 0.05fF
C4 a_159_n84# a_n129_n84# 0.05fF
C5 a_63_n84# w_n359_n303# 0.06fF
C6 a_n129_n84# a_n221_n84# 0.24fF
C7 a_n129_n84# a_n33_n84# 0.24fF
C8 a_n63_n110# a_33_n110# 0.02fF
C9 a_63_n84# a_n129_n84# 0.09fF
C10 a_129_n110# a_33_n110# 0.02fF
C11 a_159_n84# a_n221_n84# 0.04fF
C12 a_159_n84# a_n33_n84# 0.09fF
C13 a_63_n84# a_159_n84# 0.24fF
C14 a_n33_n84# a_n221_n84# 0.09fF
C15 a_n159_n110# a_n63_n110# 0.02fF
C16 a_63_n84# a_n221_n84# 0.05fF
C17 a_63_n84# a_n33_n84# 0.24fF
C18 a_159_n84# VSUBS 0.03fF
C19 a_63_n84# VSUBS 0.03fF
C20 a_n33_n84# VSUBS 0.03fF
C21 a_n129_n84# VSUBS 0.03fF
C22 a_n221_n84# VSUBS 0.03fF
C23 a_129_n110# VSUBS 0.05fF
C24 a_33_n110# VSUBS 0.05fF
C25 a_n63_n110# VSUBS 0.05fF
C26 a_n159_n110# VSUBS 0.05fF
C27 w_n359_n303# VSUBS 2.19fF
.ends

.subckt sky130_fd_pr__nfet_01v8_DXA56D w_n359_n252# a_n33_n42# a_129_n68# a_n159_n68#
+ a_n221_n42# a_159_n42# a_n129_n42# a_33_n68# a_n63_n68# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n129_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_159_n42# a_129_n68# a_63_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_n129_n42# a_n159_n68# a_n221_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n33_n42# a_159_n42# 0.05fF
C1 a_n221_n42# a_n129_n42# 0.12fF
C2 a_n33_n42# a_63_n42# 0.12fF
C3 a_n221_n42# a_n33_n42# 0.05fF
C4 a_33_n68# a_n63_n68# 0.02fF
C5 a_n129_n42# a_n33_n42# 0.12fF
C6 a_159_n42# a_63_n42# 0.12fF
C7 a_129_n68# a_33_n68# 0.02fF
C8 a_n221_n42# a_159_n42# 0.02fF
C9 a_n129_n42# a_159_n42# 0.03fF
C10 a_n159_n68# a_n63_n68# 0.02fF
C11 a_n221_n42# a_63_n42# 0.03fF
C12 a_n129_n42# a_63_n42# 0.05fF
C13 a_159_n42# w_n359_n252# 0.07fF
C14 a_63_n42# w_n359_n252# 0.06fF
C15 a_n33_n42# w_n359_n252# 0.06fF
C16 a_n129_n42# w_n359_n252# 0.06fF
C17 a_n221_n42# w_n359_n252# 0.07fF
C18 a_129_n68# w_n359_n252# 0.05fF
C19 a_33_n68# w_n359_n252# 0.05fF
C20 a_n63_n68# w_n359_n252# 0.05fF
C21 a_n159_n68# w_n359_n252# 0.05fF
.ends

.subckt inverter_min_x4 vdd in vss out
Xsky130_fd_pr__pfet_01v8_ZP3U9B_0 vss out out vdd in vdd in in vdd in out sky130_fd_pr__pfet_01v8_ZP3U9B
Xsky130_fd_pr__nfet_01v8_DXA56D_0 vss out in in out out vss in in vss sky130_fd_pr__nfet_01v8_DXA56D
C0 in vdd 0.33fF
C1 out vdd 0.62fF
C2 in out 0.67fF
C3 out vss 0.66fF
C4 in vss 1.89fF
C5 vdd vss 3.87fF
.ends

.subckt sky130_fd_pr__pfet_01v8_BDRUME VSUBS a_351_n84# a_n513_n84# a_639_n84# a_159_n84#
+ a_n321_n84# a_447_n84# a_n753_n181# a_n609_n84# w_n935_n303# a_n129_n84# a_735_n84#
+ a_255_n84# a_n417_n84# a_63_n84# a_543_n84# a_n705_n84# a_n225_n84# a_n797_n84#
+ a_n33_n84#
X0 a_n705_n84# a_n753_n181# a_n797_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_n513_n84# a_n753_n181# a_n609_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_n417_n84# a_n753_n181# a_n513_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_n321_n84# a_n753_n181# a_n417_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_n225_n84# a_n753_n181# a_n321_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 a_n129_n84# a_n753_n181# a_n225_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 a_n609_n84# a_n753_n181# a_n705_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_63_n84# a_n753_n181# a_n33_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_n33_n84# a_n753_n181# a_n129_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_159_n84# a_n753_n181# a_63_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_255_n84# a_n753_n181# a_159_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 a_351_n84# a_n753_n181# a_255_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 a_543_n84# a_n753_n181# a_447_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 a_447_n84# a_n753_n181# a_351_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 a_639_n84# a_n753_n181# a_543_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_735_n84# a_n753_n181# a_639_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_543_n84# a_255_n84# 0.05fF
C1 a_n417_n84# a_n225_n84# 0.09fF
C2 a_639_n84# a_351_n84# 0.05fF
C3 a_351_n84# a_63_n84# 0.05fF
C4 a_63_n84# a_n129_n84# 0.09fF
C5 a_543_n84# w_n935_n303# 0.03fF
C6 a_735_n84# a_447_n84# 0.05fF
C7 a_n417_n84# a_n705_n84# 0.05fF
C8 a_639_n84# a_543_n84# 0.24fF
C9 a_n417_n84# a_n797_n84# 0.04fF
C10 a_159_n84# a_351_n84# 0.09fF
C11 a_159_n84# a_n129_n84# 0.05fF
C12 a_n225_n84# a_n321_n84# 0.24fF
C13 a_n417_n84# a_n513_n84# 0.24fF
C14 a_159_n84# a_543_n84# 0.04fF
C15 a_n705_n84# a_n321_n84# 0.04fF
C16 a_n417_n84# a_n33_n84# 0.04fF
C17 a_63_n84# a_n225_n84# 0.05fF
C18 a_351_n84# a_543_n84# 0.09fF
C19 a_n705_n84# w_n935_n303# 0.04fF
C20 a_n513_n84# a_n321_n84# 0.09fF
C21 a_n797_n84# w_n935_n303# 0.08fF
C22 a_255_n84# a_447_n84# 0.09fF
C23 a_159_n84# a_n225_n84# 0.04fF
C24 a_447_n84# w_n935_n303# 0.02fF
C25 a_n513_n84# w_n935_n303# 0.02fF
C26 a_n33_n84# a_n321_n84# 0.05fF
C27 a_639_n84# a_447_n84# 0.09fF
C28 a_255_n84# a_n33_n84# 0.05fF
C29 a_n225_n84# a_n609_n84# 0.04fF
C30 a_735_n84# w_n935_n303# 0.08fF
C31 a_63_n84# a_447_n84# 0.04fF
C32 a_n225_n84# a_n129_n84# 0.24fF
C33 a_n417_n84# a_n321_n84# 0.24fF
C34 a_735_n84# a_639_n84# 0.24fF
C35 a_n609_n84# a_n705_n84# 0.24fF
C36 a_159_n84# a_447_n84# 0.05fF
C37 a_n797_n84# a_n609_n84# 0.09fF
C38 a_63_n84# a_n33_n84# 0.24fF
C39 a_n609_n84# a_n513_n84# 0.24fF
C40 a_351_n84# a_447_n84# 0.24fF
C41 a_159_n84# a_n33_n84# 0.09fF
C42 a_n129_n84# a_n513_n84# 0.04fF
C43 a_735_n84# a_351_n84# 0.04fF
C44 a_543_n84# a_447_n84# 0.24fF
C45 a_351_n84# a_n33_n84# 0.04fF
C46 a_n129_n84# a_n33_n84# 0.24fF
C47 a_63_n84# a_n321_n84# 0.04fF
C48 a_639_n84# a_255_n84# 0.04fF
C49 a_735_n84# a_543_n84# 0.09fF
C50 a_255_n84# a_63_n84# 0.09fF
C51 a_n417_n84# a_n609_n84# 0.09fF
C52 a_n417_n84# a_n129_n84# 0.05fF
C53 a_639_n84# w_n935_n303# 0.04fF
C54 a_159_n84# a_255_n84# 0.24fF
C55 a_n609_n84# a_n321_n84# 0.05fF
C56 a_n797_n84# a_n705_n84# 0.24fF
C57 a_n225_n84# a_n513_n84# 0.05fF
C58 a_n129_n84# a_n321_n84# 0.09fF
C59 a_351_n84# a_255_n84# 0.24fF
C60 a_255_n84# a_n129_n84# 0.04fF
C61 a_n705_n84# a_n513_n84# 0.09fF
C62 a_159_n84# a_63_n84# 0.24fF
C63 a_n609_n84# w_n935_n303# 0.03fF
C64 a_n225_n84# a_n33_n84# 0.09fF
C65 a_n797_n84# a_n513_n84# 0.05fF
C66 a_735_n84# VSUBS 0.03fF
C67 a_639_n84# VSUBS 0.03fF
C68 a_543_n84# VSUBS 0.03fF
C69 a_447_n84# VSUBS 0.03fF
C70 a_351_n84# VSUBS 0.03fF
C71 a_255_n84# VSUBS 0.03fF
C72 a_159_n84# VSUBS 0.03fF
C73 a_63_n84# VSUBS 0.03fF
C74 a_n33_n84# VSUBS 0.03fF
C75 a_n129_n84# VSUBS 0.03fF
C76 a_n225_n84# VSUBS 0.03fF
C77 a_n321_n84# VSUBS 0.03fF
C78 a_n417_n84# VSUBS 0.03fF
C79 a_n513_n84# VSUBS 0.03fF
C80 a_n609_n84# VSUBS 0.03fF
C81 a_n705_n84# VSUBS 0.03fF
C82 a_n797_n84# VSUBS 0.03fF
C83 a_n753_n181# VSUBS 2.56fF
C84 w_n935_n303# VSUBS 4.96fF
.ends

.subckt sky130_fd_pr__nfet_01v8_QQE8KM a_543_n42# a_n705_n42# a_n225_n42# a_n797_n42#
+ a_n33_n42# a_351_n42# a_n513_n42# a_639_n42# a_159_n42# w_n935_n252# a_n757_64#
+ a_n321_n42# a_447_n42# a_n609_n42# a_n129_n42# a_735_n42# a_255_n42# a_n417_n42#
+ a_63_n42#
X0 a_63_n42# a_n757_64# a_n33_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n757_64# a_n129_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_351_n42# a_n757_64# a_255_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_159_n42# a_n757_64# a_63_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_255_n42# a_n757_64# a_159_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_447_n42# a_n757_64# a_351_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_543_n42# a_n757_64# a_447_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_735_n42# a_n757_64# a_639_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_639_n42# a_n757_64# a_543_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_n321_n42# a_n757_64# a_n417_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_n705_n42# a_n757_64# a_n797_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_n513_n42# a_n757_64# a_n609_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_n417_n42# a_n757_64# a_n513_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_n225_n42# a_n757_64# a_n321_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_n129_n42# a_n757_64# a_n225_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_n609_n42# a_n757_64# a_n705_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_255_n42# a_543_n42# 0.03fF
C1 a_351_n42# a_447_n42# 0.12fF
C2 a_n225_n42# a_n321_n42# 0.12fF
C3 a_159_n42# a_255_n42# 0.12fF
C4 a_n129_n42# a_159_n42# 0.03fF
C5 a_447_n42# a_543_n42# 0.12fF
C6 a_639_n42# a_255_n42# 0.02fF
C7 a_n321_n42# a_n33_n42# 0.03fF
C8 a_159_n42# a_447_n42# 0.03fF
C9 a_n129_n42# a_255_n42# 0.02fF
C10 a_n417_n42# a_n321_n42# 0.12fF
C11 a_n225_n42# a_63_n42# 0.03fF
C12 a_639_n42# a_447_n42# 0.05fF
C13 a_255_n42# a_447_n42# 0.05fF
C14 a_63_n42# a_n33_n42# 0.12fF
C15 a_n513_n42# a_n321_n42# 0.05fF
C16 a_n705_n42# a_n417_n42# 0.03fF
C17 a_n321_n42# a_n609_n42# 0.03fF
C18 a_n225_n42# a_n33_n42# 0.05fF
C19 a_n417_n42# a_n225_n42# 0.05fF
C20 a_n705_n42# a_n513_n42# 0.05fF
C21 a_351_n42# a_63_n42# 0.03fF
C22 a_n417_n42# a_n33_n42# 0.02fF
C23 a_n129_n42# a_n321_n42# 0.05fF
C24 a_n513_n42# a_n225_n42# 0.03fF
C25 a_159_n42# a_63_n42# 0.12fF
C26 a_n705_n42# a_n797_n42# 0.12fF
C27 a_n705_n42# a_n609_n42# 0.12fF
C28 a_255_n42# a_63_n42# 0.05fF
C29 a_n129_n42# a_63_n42# 0.05fF
C30 a_n417_n42# a_n513_n42# 0.12fF
C31 a_n225_n42# a_n609_n42# 0.02fF
C32 a_447_n42# a_63_n42# 0.02fF
C33 a_351_n42# a_n33_n42# 0.02fF
C34 a_159_n42# a_n225_n42# 0.02fF
C35 a_n417_n42# a_n797_n42# 0.02fF
C36 a_n417_n42# a_n609_n42# 0.05fF
C37 a_159_n42# a_n33_n42# 0.05fF
C38 a_n129_n42# a_n225_n42# 0.12fF
C39 a_351_n42# a_735_n42# 0.02fF
C40 a_n797_n42# a_n513_n42# 0.03fF
C41 a_n513_n42# a_n609_n42# 0.12fF
C42 a_255_n42# a_n33_n42# 0.03fF
C43 a_n129_n42# a_n33_n42# 0.12fF
C44 a_735_n42# a_543_n42# 0.05fF
C45 a_n129_n42# a_n417_n42# 0.03fF
C46 a_639_n42# a_735_n42# 0.12fF
C47 a_351_n42# a_543_n42# 0.05fF
C48 a_n797_n42# a_n609_n42# 0.05fF
C49 a_63_n42# a_n321_n42# 0.02fF
C50 a_n129_n42# a_n513_n42# 0.02fF
C51 a_351_n42# a_159_n42# 0.05fF
C52 a_351_n42# a_639_n42# 0.03fF
C53 a_159_n42# a_543_n42# 0.02fF
C54 a_447_n42# a_735_n42# 0.03fF
C55 a_n705_n42# a_n321_n42# 0.02fF
C56 a_351_n42# a_255_n42# 0.12fF
C57 a_639_n42# a_543_n42# 0.12fF
C58 a_735_n42# w_n935_n252# 0.07fF
C59 a_639_n42# w_n935_n252# 0.05fF
C60 a_543_n42# w_n935_n252# 0.05fF
C61 a_447_n42# w_n935_n252# 0.04fF
C62 a_351_n42# w_n935_n252# 0.04fF
C63 a_255_n42# w_n935_n252# 0.04fF
C64 a_159_n42# w_n935_n252# 0.04fF
C65 a_63_n42# w_n935_n252# 0.04fF
C66 a_n33_n42# w_n935_n252# 0.04fF
C67 a_n129_n42# w_n935_n252# 0.04fF
C68 a_n225_n42# w_n935_n252# 0.04fF
C69 a_n321_n42# w_n935_n252# 0.04fF
C70 a_n417_n42# w_n935_n252# 0.04fF
C71 a_n513_n42# w_n935_n252# 0.04fF
C72 a_n609_n42# w_n935_n252# 0.05fF
C73 a_n705_n42# w_n935_n252# 0.05fF
C74 a_n797_n42# w_n935_n252# 0.07fF
C75 a_n757_64# w_n935_n252# 2.44fF
.ends

.subckt inverter_min_x16 in out vss vdd
Xsky130_fd_pr__pfet_01v8_BDRUME_0 vss out vdd vdd out vdd vdd in out vdd vdd out vdd
+ out vdd out vdd out out out sky130_fd_pr__pfet_01v8_BDRUME
Xsky130_fd_pr__nfet_01v8_QQE8KM_0 out vss out out out out vss vss out vss in vss vss
+ out vss out vss out vss sky130_fd_pr__nfet_01v8_QQE8KM
C0 in out 1.40fF
C1 vdd out 1.63fF
C2 vdd in 1.15fF
C3 out vss 0.98fF
C4 in vss 7.30fF
C5 vdd vss 10.49fF
.ends

.subckt sky130_fd_pr__pfet_01v8_75PKJG VSUBS a_n33_n102# w_n359_n321# a_n177_n199#
+ a_63_n102# a_n129_n102# a_n221_n102# a_25_n199# a_159_n102#
X0 a_159_n102# a_25_n199# a_63_n102# w_n359_n321# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
X1 a_63_n102# a_25_n199# a_n33_n102# w_n359_n321# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
X2 a_n129_n102# a_n177_n199# a_n221_n102# w_n359_n321# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
X3 a_n33_n102# a_n177_n199# a_n129_n102# w_n359_n321# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
C0 a_63_n102# a_159_n102# 0.30fF
C1 a_63_n102# a_n221_n102# 0.07fF
C2 a_n33_n102# a_n129_n102# 0.30fF
C3 w_n359_n321# a_n129_n102# 0.07fF
C4 a_n177_n199# a_25_n199# 0.07fF
C5 a_159_n102# a_n129_n102# 0.07fF
C6 a_n221_n102# a_n129_n102# 0.30fF
C7 a_63_n102# a_n129_n102# 0.11fF
C8 a_n33_n102# w_n359_n321# 0.06fF
C9 a_n33_n102# a_159_n102# 0.11fF
C10 a_n221_n102# a_n33_n102# 0.11fF
C11 w_n359_n321# a_159_n102# 0.10fF
C12 a_n221_n102# w_n359_n321# 0.10fF
C13 a_n221_n102# a_159_n102# 0.05fF
C14 a_63_n102# a_n33_n102# 0.30fF
C15 a_63_n102# w_n359_n321# 0.07fF
C16 a_159_n102# VSUBS 0.03fF
C17 a_63_n102# VSUBS 0.03fF
C18 a_n33_n102# VSUBS 0.03fF
C19 a_n129_n102# VSUBS 0.03fF
C20 a_n221_n102# VSUBS 0.03fF
C21 a_25_n199# VSUBS 0.22fF
C22 a_n177_n199# VSUBS 0.22fF
C23 w_n359_n321# VSUBS 2.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_XRJ78J a_n33_n102# w_n263_n312# a_63_n102# a_n125_n102#
+ a_n81_124#
X0 a_n33_n102# a_n81_124# a_n125_n102# w_n263_n312# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
X1 a_63_n102# a_n81_124# a_n33_n102# w_n263_n312# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
C0 a_63_n102# a_n125_n102# 0.11fF
C1 a_n33_n102# a_n125_n102# 0.30fF
C2 a_n33_n102# a_63_n102# 0.30fF
C3 a_63_n102# w_n263_n312# 0.06fF
C4 a_n33_n102# w_n263_n312# 0.08fF
C5 a_n125_n102# w_n263_n312# 0.12fF
C6 a_n81_124# w_n263_n312# 0.21fF
.ends

.subckt nand_logic avss1p8 in1 avdd1p8 in2 out m1_21_n341#
Xsky130_fd_pr__pfet_01v8_75PKJG_0 avss1p8 avdd1p8 avdd1p8 in1 out out avdd1p8 in2
+ avdd1p8 sky130_fd_pr__pfet_01v8_75PKJG
Xsky130_fd_pr__nfet_01v8_XRJ78J_0 m1_21_n341# avss1p8 avss1p8 avss1p8 in1 sky130_fd_pr__nfet_01v8_XRJ78J
Xsky130_fd_pr__nfet_01v8_XRJ78J_1 out avss1p8 m1_21_n341# m1_21_n341# in2 sky130_fd_pr__nfet_01v8_XRJ78J
C0 avdd1p8 out 0.20fF
C1 in1 out 0.10fF
C2 in2 avdd1p8 0.02fF
C3 in2 out 0.37fF
C4 m1_21_n341# avdd1p8 0.01fF
C5 m1_21_n341# out 0.13fF
C6 in2 in1 0.07fF
C7 m1_21_n341# in1 0.25fF
C8 m1_21_n341# avss1p8 0.92fF
C9 out avss1p8 0.47fF
C10 in2 avss1p8 0.91fF
C11 in1 avss1p8 0.93fF
C12 avdd1p8 avss1p8 2.37fF
.ends

.subckt res_amp_sync_v2 avdd1p8 DFlipFlop_4/Q vss clkn DFlipFlop_4/latch_diff_1/m1_657_280#
+ DFlipFlop_4/nQ DFlipFlop_3/latch_diff_1/nD DFlipFlop_3/latch_diff_0/D DFlipFlop_3/Q
+ DFlipFlop_3/D DFlipFlop_4/D DFlipFlop_1/D DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_4/latch_diff_1/D DFlipFlop_4/latch_diff_1/nD DFlipFlop_4/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_4/latch_diff_0/D DFlipFlop_3/latch_diff_1/D clk_amp DFlipFlop_3/nQ clkp
+ rst
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vss avdd1p8 DFlipFlop_0/latch_diff_1/D
+ DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_0/nQ clkn DFlipFlop_0/latch_diff_0/nD
+ DFlipFlop_0/Q DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/latch_diff_1/m1_657_280# DFlipFlop_3/D
+ DFlipFlop_0/latch_diff_0/D clkp DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_1 DFlipFlop_1/latch_diff_0/m1_657_280# vss avdd1p8 DFlipFlop_1/latch_diff_1/D
+ DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_1/nQ DFlipFlop_0/Q DFlipFlop_1/latch_diff_0/nD
+ DFlipFlop_2/D DFlipFlop_1/latch_diff_1/nD DFlipFlop_1/latch_diff_1/m1_657_280# DFlipFlop_1/D
+ DFlipFlop_1/latch_diff_0/D DFlipFlop_3/D DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_2 DFlipFlop_2/latch_diff_0/m1_657_280# vss avdd1p8 DFlipFlop_2/latch_diff_1/D
+ DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_2/nQ clkn DFlipFlop_2/latch_diff_0/nD
+ DFlipFlop_2/Q DFlipFlop_2/latch_diff_1/nD DFlipFlop_2/latch_diff_1/m1_657_280# DFlipFlop_2/D
+ DFlipFlop_2/latch_diff_0/D clkp DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_3 DFlipFlop_3/latch_diff_0/m1_657_280# vss avdd1p8 DFlipFlop_3/latch_diff_1/D
+ DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_3/nQ clkn DFlipFlop_3/latch_diff_0/nD
+ DFlipFlop_3/Q DFlipFlop_3/latch_diff_1/nD DFlipFlop_3/latch_diff_1/m1_657_280# DFlipFlop_3/D
+ DFlipFlop_3/latch_diff_0/D clkp DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
Xinverter_min_x4_0 avdd1p8 DFlipFlop_0/Q vss DFlipFlop_3/D inverter_min_x4
Xinverter_min_x4_1 avdd1p8 nand_logic_0/out vss DFlipFlop_4/D inverter_min_x4
XDFlipFlop_4 DFlipFlop_4/latch_diff_0/m1_657_280# vss avdd1p8 DFlipFlop_4/latch_diff_1/D
+ DFlipFlop_4/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_4/nQ clkn DFlipFlop_4/latch_diff_0/nD
+ DFlipFlop_4/Q DFlipFlop_4/latch_diff_1/nD DFlipFlop_4/latch_diff_1/m1_657_280# DFlipFlop_4/D
+ DFlipFlop_4/latch_diff_0/D clkp DFlipFlop_4/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
Xinverter_min_x4_2 avdd1p8 DFlipFlop_2/D vss DFlipFlop_1/D inverter_min_x4
Xinverter_min_x4_3 avdd1p8 nand_logic_1/out vss rst inverter_min_x4
Xinverter_min_x4_4 avdd1p8 DFlipFlop_4/Q vss inverter_min_x4_4/out inverter_min_x4
Xinverter_min_x16_0 inverter_min_x4_4/out clk_amp vss avdd1p8 inverter_min_x16
Xnand_logic_0 vss DFlipFlop_2/Q avdd1p8 DFlipFlop_3/Q nand_logic_0/out nand_logic_0/m1_21_n341#
+ nand_logic
Xnand_logic_1 vss DFlipFlop_4/D avdd1p8 clkp nand_logic_1/out nand_logic_1/m1_21_n341#
+ nand_logic
C0 clkp nand_logic_1/out 0.03fF
C1 DFlipFlop_3/nQ avdd1p8 0.03fF
C2 clkp DFlipFlop_2/nQ 0.13fF
C3 DFlipFlop_1/latch_diff_0/m1_657_280# DFlipFlop_3/D 0.28fF
C4 DFlipFlop_3/D DFlipFlop_2/D 0.06fF
C5 DFlipFlop_3/D DFlipFlop_0/latch_diff_1/D 0.08fF
C6 DFlipFlop_1/D DFlipFlop_1/nQ 0.02fF
C7 DFlipFlop_3/Q DFlipFlop_2/nQ 0.02fF
C8 clkn DFlipFlop_4/nQ 0.02fF
C9 clkn DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in 0.14fF
C10 DFlipFlop_0/Q avdd1p8 0.66fF
C11 DFlipFlop_2/latch_diff_0/D DFlipFlop_2/D -0.07fF
C12 clkn DFlipFlop_3/latch_diff_1/nD 0.17fF
C13 nand_logic_1/out DFlipFlop_4/D 0.01fF
C14 clkp DFlipFlop_4/latch_diff_0/m1_657_280# 0.30fF
C15 DFlipFlop_2/D avdd1p8 4.16fF
C16 clkp DFlipFlop_0/latch_diff_0/nD 0.08fF
C17 nand_logic_0/out DFlipFlop_2/Q 0.02fF
C18 clkn DFlipFlop_3/D 0.35fF
C19 DFlipFlop_3/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.43fF
C20 clkn DFlipFlop_4/clock_inverter_0/inverter_cp_x1_2/in -0.33fF
C21 nand_logic_0/out avdd1p8 0.03fF
C22 DFlipFlop_1/latch_diff_1/D DFlipFlop_0/Q 0.10fF
C23 avdd1p8 clk_amp 0.10fF
C24 clkn DFlipFlop_4/latch_diff_1/D 0.08fF
C25 clkp DFlipFlop_3/Q 0.17fF
C26 DFlipFlop_0/latch_diff_0/D DFlipFlop_3/D 0.31fF
C27 clkp DFlipFlop_3/latch_diff_0/m1_657_280# 0.30fF
C28 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_0/Q 0.55fF
C29 clkn DFlipFlop_0/nQ 0.02fF
C30 clkn DFlipFlop_2/latch_diff_0/D 0.12fF
C31 nand_logic_0/m1_21_n341# DFlipFlop_3/Q 0.07fF
C32 clkp DFlipFlop_2/latch_diff_0/m1_657_280# 0.30fF
C33 DFlipFlop_4/latch_diff_1/nD clkn 0.17fF
C34 clkp DFlipFlop_4/D 0.24fF
C35 inverter_min_x4_4/out avdd1p8 0.09fF
C36 clkn avdd1p8 -1.00fF
C37 avdd1p8 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.01fF
C38 DFlipFlop_0/Q DFlipFlop_1/latch_diff_1/nD 0.19fF
C39 nand_logic_0/m1_21_n341# DFlipFlop_4/D 0.02fF
C40 clkn DFlipFlop_3/latch_diff_1/D 0.08fF
C41 DFlipFlop_4/Q inverter_min_x4_4/out 0.01fF
C42 DFlipFlop_3/Q DFlipFlop_4/D 0.94fF
C43 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_2/D 0.49fF
C44 clkp DFlipFlop_4/latch_diff_0/nD 0.08fF
C45 clkn DFlipFlop_0/latch_diff_1/nD 0.17fF
C46 clkp DFlipFlop_4/nQ 0.02fF
C47 DFlipFlop_1/D DFlipFlop_3/D 0.28fF
C48 clkn DFlipFlop_3/nQ 0.10fF
C49 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out avdd1p8 0.01fF
C50 clkp DFlipFlop_3/latch_diff_1/nD 0.10fF
C51 clkn DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in 0.14fF
C52 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out avdd1p8 0.01fF
C53 nand_logic_1/out avdd1p8 0.04fF
C54 clkp DFlipFlop_3/D 0.35fF
C55 DFlipFlop_1/nQ DFlipFlop_3/D 0.05fF
C56 rst avdd1p8 0.02fF
C57 clkp DFlipFlop_4/latch_diff_1/D 0.15fF
C58 DFlipFlop_1/D avdd1p8 2.55fF
C59 clkn DFlipFlop_4/latch_diff_1/m1_657_280# 0.30fF
C60 clkp DFlipFlop_0/nQ 0.02fF
C61 DFlipFlop_2/latch_diff_1/D DFlipFlop_2/D 0.03fF
C62 DFlipFlop_3/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.54fF
C63 clkp DFlipFlop_4/latch_diff_1/nD 0.10fF
C64 clkn DFlipFlop_2/D 0.15fF
C65 clkn DFlipFlop_0/latch_diff_1/D 0.08fF
C66 inverter_min_x4_4/out clk_amp 0.12fF
C67 clkp DFlipFlop_2/Q 0.11fF
C68 clkp avdd1p8 0.53fF
C69 DFlipFlop_1/D DFlipFlop_1/latch_diff_1/D 0.02fF
C70 clkn DFlipFlop_4/latch_diff_0/D 0.12fF
C71 clkp DFlipFlop_3/latch_diff_1/D 0.15fF
C72 DFlipFlop_1/D DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in 0.41fF
C73 clkp DFlipFlop_4/Q 0.20fF
C74 DFlipFlop_2/latch_diff_1/nD clkn 0.17fF
C75 DFlipFlop_1/latch_diff_0/D DFlipFlop_0/Q 0.74fF
C76 DFlipFlop_3/Q DFlipFlop_2/Q 0.09fF
C77 DFlipFlop_3/Q avdd1p8 0.76fF
C78 clkn DFlipFlop_2/latch_diff_1/D 0.08fF
C79 clkp DFlipFlop_0/latch_diff_1/nD 0.10fF
C80 clkp DFlipFlop_2/latch_diff_0/nD 0.08fF
C81 nand_logic_1/out nand_logic_1/m1_21_n341# 0.01fF
C82 DFlipFlop_3/Q DFlipFlop_4/Q 0.11fF
C83 clkp DFlipFlop_4/clock_inverter_0/inverter_cp_x1_0/out -0.31fF
C84 clkn DFlipFlop_0/latch_diff_0/D 0.12fF
C85 rst nand_logic_1/m1_21_n341# 0.02fF
C86 DFlipFlop_4/D avdd1p8 0.52fF
C87 clkn DFlipFlop_3/latch_diff_1/m1_657_280# 0.30fF
C88 clkp DFlipFlop_3/nQ 0.13fF
C89 DFlipFlop_1/D DFlipFlop_0/Q 0.72fF
C90 DFlipFlop_4/Q DFlipFlop_4/D 0.27fF
C91 DFlipFlop_2/D DFlipFlop_2/nQ 0.03fF
C92 DFlipFlop_1/latch_diff_1/m1_657_280# DFlipFlop_0/Q 0.25fF
C93 clkn DFlipFlop_2/latch_diff_1/m1_657_280# 0.30fF
C94 DFlipFlop_1/D DFlipFlop_2/D 0.02fF
C95 clkp nand_logic_1/m1_21_n341# 0.09fF
C96 DFlipFlop_1/nQ DFlipFlop_0/Q 0.01fF
C97 clkp DFlipFlop_0/latch_diff_0/m1_657_280# 0.32fF
C98 DFlipFlop_4/D DFlipFlop_4/clock_inverter_0/inverter_cp_x1_0/out 0.42fF
C99 clkn DFlipFlop_2/nQ 0.02fF
C100 clkp DFlipFlop_2/D 0.15fF
C101 clkp DFlipFlop_0/latch_diff_1/D 0.15fF
C102 DFlipFlop_0/nQ DFlipFlop_3/D 0.08fF
C103 clkp clk_amp 0.52fF
C104 DFlipFlop_4/nQ DFlipFlop_4/Q 0.06fF
C105 nand_logic_0/out nand_logic_0/m1_21_n341# 0.01fF
C106 DFlipFlop_4/D nand_logic_1/m1_21_n341# 0.09fF
C107 DFlipFlop_3/D avdd1p8 4.16fF
C108 DFlipFlop_4/clock_inverter_0/inverter_cp_x1_2/in avdd1p8 0.03fF
C109 nand_logic_0/out DFlipFlop_3/Q 0.01fF
C110 DFlipFlop_2/latch_diff_1/nD clkp 0.20fF
C111 clkp DFlipFlop_2/latch_diff_1/D 0.15fF
C112 clkp inverter_min_x4_4/out 0.43fF
C113 DFlipFlop_3/latch_diff_0/nD clkp 0.08fF
C114 clkp clkn 0.22fF
C115 clkp DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.16fF
C116 nand_logic_0/out DFlipFlop_4/D 0.04fF
C117 DFlipFlop_0/latch_diff_1/nD DFlipFlop_3/D 0.17fF
C118 DFlipFlop_3/Q DFlipFlop_2/latch_diff_1/D 0.03fF
C119 DFlipFlop_1/latch_diff_1/D DFlipFlop_3/D 0.03fF
C120 clkn DFlipFlop_3/latch_diff_0/D 0.12fF
C121 DFlipFlop_2/Q avdd1p8 0.05fF
C122 clkn DFlipFlop_3/Q 0.12fF
C123 clkn DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.14fF
C124 DFlipFlop_4/Q avdd1p8 4.03fF
C125 nand_logic_1/out rst 0.04fF
C126 DFlipFlop_0/latch_diff_1/m1_657_280# clkn 0.30fF
C127 clkn DFlipFlop_4/D 0.15fF
C128 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out clkp 0.16fF
C129 DFlipFlop_3/D DFlipFlop_1/latch_diff_1/nD 0.02fF
C130 DFlipFlop_0/Q DFlipFlop_3/D 0.38fF
C131 avdd1p8 DFlipFlop_4/clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C132 clkp DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out 0.16fF
C133 DFlipFlop_3/Q DFlipFlop_2/latch_diff_1/m1_657_280# 0.04fF
C134 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in avdd1p8 0.02fF
C135 nand_logic_1/m1_21_n341# vss 0.86fF
C136 nand_logic_0/m1_21_n341# vss 0.90fF
C137 clk_amp vss 0.43fF
C138 inverter_min_x4_4/out vss 5.90fF
C139 rst vss 0.71fF
C140 nand_logic_1/out vss 1.76fF
C141 DFlipFlop_4/Q vss -2.08fF
C142 DFlipFlop_4/latch_diff_1/m1_657_280# vss 0.57fF
C143 DFlipFlop_4/nQ vss 0.48fF
C144 DFlipFlop_4/latch_diff_1/D vss -1.73fF
C145 DFlipFlop_4/latch_diff_0/m1_657_280# vss 0.57fF
C146 DFlipFlop_4/latch_diff_1/nD vss 0.57fF
C147 DFlipFlop_4/clock_inverter_0/inverter_cp_x1_2/in vss 1.94fF
C148 DFlipFlop_4/latch_diff_0/D vss 0.96fF
C149 DFlipFlop_4/clock_inverter_0/inverter_cp_x1_0/out vss 1.84fF
C150 DFlipFlop_4/D vss 4.59fF
C151 DFlipFlop_4/latch_diff_0/nD vss 1.14fF
C152 nand_logic_0/out vss 1.26fF
C153 DFlipFlop_3/Q vss -2.01fF
C154 DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.72fF
C155 clkn vss -2.25fF
C156 DFlipFlop_3/nQ vss 0.50fF
C157 DFlipFlop_3/latch_diff_1/D vss -1.72fF
C158 DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C159 clkp vss -22.80fF
C160 DFlipFlop_3/latch_diff_1/nD vss 0.58fF
C161 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C162 DFlipFlop_3/latch_diff_0/D vss 0.96fF
C163 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C164 DFlipFlop_3/D vss 1.64fF
C165 avdd1p8 vss 196.01fF
C166 DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C167 DFlipFlop_2/Q vss -1.05fF
C168 DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.65fF
C169 DFlipFlop_2/nQ vss 0.48fF
C170 DFlipFlop_2/latch_diff_1/D vss -1.73fF
C171 DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C172 DFlipFlop_2/latch_diff_1/nD vss 0.58fF
C173 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C174 DFlipFlop_2/latch_diff_0/D vss 0.96fF
C175 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C176 DFlipFlop_2/D vss -0.35fF
C177 DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C178 DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.59fF
C179 DFlipFlop_1/nQ vss 0.48fF
C180 DFlipFlop_1/latch_diff_1/D vss -1.73fF
C181 DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C182 DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C183 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.89fF
C184 DFlipFlop_1/latch_diff_0/D vss 0.96fF
C185 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C186 DFlipFlop_1/D vss -1.00fF
C187 DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C188 DFlipFlop_0/Q vss -3.86fF
C189 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.59fF
C190 DFlipFlop_0/nQ vss 0.48fF
C191 DFlipFlop_0/latch_diff_1/D vss -1.73fF
C192 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C193 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C194 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C195 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C196 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C197 DFlipFlop_0/latch_diff_0/nD vss 1.14fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_4L9VGG VSUBS a_291_n200# w_n487_n419# a_35_n200#
+ a_n291_n238# a_n93_n200# a_163_n200# a_n349_n200# a_n221_n200#
X0 a_291_n200# a_n291_n238# a_163_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X1 a_n221_n200# a_n291_n238# a_n349_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X2 a_35_n200# a_n291_n238# a_n93_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X3 a_163_n200# a_n291_n238# a_35_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X4 a_n93_n200# a_n291_n238# a_n221_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
C0 a_n93_n200# a_n291_n238# 0.08fF
C1 a_n349_n200# a_35_n200# 0.09fF
C2 a_n349_n200# a_n221_n200# 0.36fF
C3 a_n349_n200# w_n487_n419# 0.18fF
C4 a_n93_n200# a_n349_n200# 0.15fF
C5 a_291_n200# a_35_n200# 0.15fF
C6 a_291_n200# a_163_n200# 0.36fF
C7 a_291_n200# w_n487_n419# 0.18fF
C8 a_n93_n200# a_291_n200# 0.09fF
C9 a_35_n200# a_163_n200# 0.36fF
C10 a_n221_n200# a_35_n200# 0.15fF
C11 a_35_n200# w_n487_n419# 0.06fF
C12 a_35_n200# a_n291_n238# 0.08fF
C13 a_n221_n200# a_163_n200# 0.09fF
C14 a_n93_n200# a_35_n200# 0.36fF
C15 w_n487_n419# a_163_n200# 0.08fF
C16 a_n221_n200# w_n487_n419# 0.08fF
C17 a_n291_n238# a_163_n200# 0.08fF
C18 a_n93_n200# a_163_n200# 0.15fF
C19 a_n221_n200# a_n291_n238# 0.08fF
C20 a_n93_n200# a_n221_n200# 0.36fF
C21 w_n487_n419# a_n291_n238# 0.30fF
C22 a_n93_n200# w_n487_n419# 0.06fF
C23 a_291_n200# VSUBS 0.03fF
C24 a_163_n200# VSUBS 0.03fF
C25 a_35_n200# VSUBS 0.03fF
C26 a_n93_n200# VSUBS 0.03fF
C27 a_n221_n200# VSUBS 0.03fF
C28 a_n349_n200# VSUBS 0.03fF
C29 a_n291_n238# VSUBS 0.72fF
C30 w_n487_n419# VSUBS 4.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_L78GGD a_n73_n73# w_n211_n221# a_15_n73# a_n33_33#
X0 a_15_n73# a_n33_33# a_n73_n73# w_n211_n221# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n33_33# a_15_n73# 0.02fF
C1 a_n73_n73# a_15_n73# 0.15fF
C2 a_n33_33# a_n73_n73# 0.02fF
C3 a_15_n73# w_n211_n221# 0.11fF
C4 a_n73_n73# w_n211_n221# 0.11fF
C5 a_n33_33# w_n211_n221# 0.18fF
.ends

.subckt sky130_fd_pr__pfet_01v8_6RX2PQ VSUBS w_n211_n268# a_15_n48# a_n33_n145# a_n73_n48#
X0 a_15_n48# a_n33_n145# a_n73_n48# w_n211_n268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 w_n211_n268# a_15_n48# 0.13fF
C1 w_n211_n268# a_n73_n48# 0.13fF
C2 a_n33_n145# a_15_n48# 0.01fF
C3 a_n33_n145# a_n73_n48# 0.01fF
C4 w_n211_n268# a_n33_n145# 0.06fF
C5 a_n73_n48# a_15_n48# 0.29fF
C6 a_15_n48# VSUBS 0.03fF
C7 a_n73_n48# VSUBS 0.03fF
C8 a_n33_n145# VSUBS 0.12fF
C9 w_n211_n268# VSUBS 1.50fF
.ends

.subckt inverter_min vdd out in vss
XXM1 vss vss out in sky130_fd_pr__nfet_01v8_L78GGD
XXM2 vss vdd out in vdd sky130_fd_pr__pfet_01v8_6RX2PQ
C0 out vdd 0.20fF
C1 vdd in 0.13fF
C2 out in 0.67fF
C3 out vss 0.52fF
C4 in vss 0.72fF
C5 vdd vss 2.55fF
.ends

.subckt buffer_no_inv_x05 VSUBS in avdd1p8 inverter_min_1/in out
Xinverter_min_1 avdd1p8 out inverter_min_1/in VSUBS inverter_min
Xinverter_min_0 avdd1p8 inverter_min_1/in in VSUBS inverter_min
C0 inverter_min_1/in avdd1p8 0.09fF
C1 avdd1p8 out 0.02fF
C2 in inverter_min_1/in 0.07fF
C3 inverter_min_1/in out 0.12fF
C4 in VSUBS 0.63fF
C5 avdd1p8 VSUBS 4.78fF
C6 out VSUBS 0.45fF
C7 inverter_min_1/in VSUBS 1.08fF
.ends

.subckt sky130_fd_pr__pfet_01v8_XA7ZMQ VSUBS a_21_142# a_63_n111# a_n87_142# a_n125_n111#
+ w_n263_n330# a_n33_n111#
X0 a_n33_n111# a_n87_142# a_n125_n111# w_n263_n330# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.11e+06u l=150000u
X1 a_63_n111# a_21_142# a_n33_n111# w_n263_n330# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.11e+06u l=150000u
C0 a_n125_n111# a_n87_142# 0.02fF
C1 a_21_142# a_63_n111# 0.02fF
C2 a_n125_n111# a_n33_n111# 0.32fF
C3 w_n263_n330# a_21_142# 0.05fF
C4 a_n125_n111# a_63_n111# 0.12fF
C5 w_n263_n330# a_n87_142# 0.05fF
C6 a_n33_n111# a_63_n111# 0.32fF
C7 a_n125_n111# w_n263_n330# 0.14fF
C8 a_21_142# a_n87_142# 0.14fF
C9 a_n33_n111# w_n263_n330# 0.10fF
C10 w_n263_n330# a_63_n111# 0.14fF
C11 a_63_n111# VSUBS 0.03fF
C12 a_n33_n111# VSUBS 0.03fF
C13 a_n125_n111# VSUBS 0.03fF
C14 a_21_142# VSUBS 0.16fF
C15 a_n87_142# VSUBS 0.16fF
C16 w_n263_n330# VSUBS 2.11fF
.ends

.subckt sky130_fd_pr__nfet_01v8_HAN8QX a_15_n142# a_n33_102# a_n73_n142# w_n211_n290#
X0 a_15_n142# a_n33_102# a_n73_n142# w_n211_n290# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.11e+06u l=150000u
C0 a_n33_102# a_15_n142# 0.03fF
C1 a_n33_102# a_n73_n142# 0.03fF
C2 a_15_n142# a_n73_n142# 0.38fF
C3 a_15_n142# w_n211_n290# 0.19fF
C4 a_n73_n142# w_n211_n290# 0.19fF
C5 a_n33_102# w_n211_n290# 0.21fF
.ends

.subckt mux_2to1_logic sel avdd1p8 sel_b w_947_n633# avss1p8 out DinA DinB
Xinverter_min_0 avdd1p8 sel_b sel avss1p8 inverter_min
Xsky130_fd_pr__pfet_01v8_XA7ZMQ_0 avss1p8 sel DinA sel DinA avdd1p8 out sky130_fd_pr__pfet_01v8_XA7ZMQ
Xsky130_fd_pr__pfet_01v8_XA7ZMQ_1 avss1p8 sel_b DinB sel_b DinB avdd1p8 out sky130_fd_pr__pfet_01v8_XA7ZMQ
Xsky130_fd_pr__nfet_01v8_HAN8QX_0 out sel_b DinA avss1p8 sky130_fd_pr__nfet_01v8_HAN8QX
Xsky130_fd_pr__nfet_01v8_HAN8QX_1 out sel DinB avss1p8 sky130_fd_pr__nfet_01v8_HAN8QX
C0 DinB sel 0.02fF
C1 out DinA 0.30fF
C2 out avdd1p8 0.23fF
C3 sel_b DinA 0.56fF
C4 sel_b avdd1p8 0.74fF
C5 out sel 0.53fF
C6 sel_b sel 0.32fF
C7 DinA avdd1p8 0.26fF
C8 DinA sel 0.07fF
C9 avdd1p8 sel 0.72fF
C10 out DinB 0.37fF
C11 sel_b DinB 0.27fF
C12 DinA DinB 0.07fF
C13 avdd1p8 DinB 0.16fF
C14 out sel_b 0.58fF
C15 DinA avss1p8 0.63fF
C16 out avss1p8 1.11fF
C17 DinB avss1p8 -0.09fF
C18 sel_b avss1p8 2.16fF
C19 sel avss1p8 2.55fF
C20 avdd1p8 avss1p8 8.26fF
.ends

.subckt delay_cell_buff buffer_no_inv_x05_2/inverter_min_1/in reg2 avss1p8 mux_2to1_logic_4/DinA
+ avdd1p8 buffer_no_inv_x05_13/in clk mux_2to1_logic_3/DinA clk_out mux_2to1_logic_3/DinB
+ reg0 buffer_no_inv_x05_10/inverter_min_1/in reg1 buffer_no_inv_x05_7/inverter_min_1/in
+ nand_logic_0/in1 mux_2to1_logic_2/out mux_2to1_logic_4/sel_b mux_2to1_logic_4/out
+ mux_2to1_logic_1/DinA mux_2to1_logic_1/sel_b buffer_no_inv_x05_3/in mux_2to1_logic_5/out
+ mux_2to1_logic_0/out mux_2to1_logic_4/DinB mux_2to1_logic_3/out buffer_no_inv_x05_13/inverter_min_1/in
+ mux_2to1_logic_1/out mux_2to1_logic_5/w_947_n633# buffer_no_inv_x05_12/inverter_min_1/in
+ nand_logic_0/m1_21_n341#
Xbuffer_no_inv_x05_8 avss1p8 mux_2to1_logic_3/DinA avdd1p8 buffer_no_inv_x05_8/inverter_min_1/in
+ buffer_no_inv_x05_9/in buffer_no_inv_x05
Xbuffer_no_inv_x05_9 avss1p8 buffer_no_inv_x05_9/in avdd1p8 buffer_no_inv_x05_9/inverter_min_1/in
+ mux_2to1_logic_3/DinB buffer_no_inv_x05
Xmux_2to1_logic_0 reg2 avdd1p8 mux_2to1_logic_0/sel_b mux_2to1_logic_0/w_947_n633#
+ avss1p8 mux_2to1_logic_0/out clk mux_2to1_logic_0/DinB mux_2to1_logic
Xmux_2to1_logic_1 reg2 avdd1p8 mux_2to1_logic_1/sel_b mux_2to1_logic_1/w_947_n633#
+ avss1p8 mux_2to1_logic_1/out mux_2to1_logic_1/DinA mux_2to1_logic_1/DinB mux_2to1_logic
Xmux_2to1_logic_2 reg1 avdd1p8 mux_2to1_logic_2/sel_b mux_2to1_logic_2/w_947_n633#
+ avss1p8 mux_2to1_logic_2/out mux_2to1_logic_0/out mux_2to1_logic_1/out mux_2to1_logic
Xmux_2to1_logic_3 reg2 avdd1p8 mux_2to1_logic_3/sel_b mux_2to1_logic_3/w_947_n633#
+ avss1p8 mux_2to1_logic_3/out mux_2to1_logic_3/DinA mux_2to1_logic_3/DinB mux_2to1_logic
Xmux_2to1_logic_4 reg2 avdd1p8 mux_2to1_logic_4/sel_b mux_2to1_logic_4/w_947_n633#
+ avss1p8 mux_2to1_logic_4/out mux_2to1_logic_4/DinA mux_2to1_logic_4/DinB mux_2to1_logic
Xmux_2to1_logic_5 reg1 avdd1p8 mux_2to1_logic_5/sel_b mux_2to1_logic_5/w_947_n633#
+ avss1p8 mux_2to1_logic_5/out mux_2to1_logic_3/out mux_2to1_logic_4/out mux_2to1_logic
Xmux_2to1_logic_6 reg0 avdd1p8 mux_2to1_logic_6/sel_b mux_2to1_logic_6/w_947_n633#
+ avss1p8 nand_logic_0/in1 mux_2to1_logic_2/out mux_2to1_logic_5/out mux_2to1_logic
Xbuffer_no_inv_x05_10 avss1p8 mux_2to1_logic_3/DinB avdd1p8 buffer_no_inv_x05_10/inverter_min_1/in
+ buffer_no_inv_x05_11/in buffer_no_inv_x05
Xnand_logic_0 avss1p8 nand_logic_0/in1 avdd1p8 clk clk_out nand_logic_0/m1_21_n341#
+ nand_logic
Xbuffer_no_inv_x05_11 avss1p8 buffer_no_inv_x05_11/in avdd1p8 buffer_no_inv_x05_11/inverter_min_1/in
+ mux_2to1_logic_4/DinA buffer_no_inv_x05
Xbuffer_no_inv_x05_12 avss1p8 mux_2to1_logic_4/DinA avdd1p8 buffer_no_inv_x05_12/inverter_min_1/in
+ buffer_no_inv_x05_13/in buffer_no_inv_x05
Xbuffer_no_inv_x05_13 avss1p8 buffer_no_inv_x05_13/in avdd1p8 buffer_no_inv_x05_13/inverter_min_1/in
+ mux_2to1_logic_4/DinB buffer_no_inv_x05
Xbuffer_no_inv_x05_0 avss1p8 clk avdd1p8 buffer_no_inv_x05_0/inverter_min_1/in buffer_no_inv_x05_1/in
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_2 avss1p8 mux_2to1_logic_0/DinB avdd1p8 buffer_no_inv_x05_2/inverter_min_1/in
+ buffer_no_inv_x05_3/in buffer_no_inv_x05
Xbuffer_no_inv_x05_1 avss1p8 buffer_no_inv_x05_1/in avdd1p8 buffer_no_inv_x05_1/inverter_min_1/in
+ mux_2to1_logic_0/DinB buffer_no_inv_x05
Xbuffer_no_inv_x05_3 avss1p8 buffer_no_inv_x05_3/in avdd1p8 buffer_no_inv_x05_3/inverter_min_1/in
+ mux_2to1_logic_1/DinA buffer_no_inv_x05
Xbuffer_no_inv_x05_4 avss1p8 mux_2to1_logic_1/DinA avdd1p8 buffer_no_inv_x05_4/inverter_min_1/in
+ buffer_no_inv_x05_5/in buffer_no_inv_x05
Xbuffer_no_inv_x05_5 avss1p8 buffer_no_inv_x05_5/in avdd1p8 buffer_no_inv_x05_5/inverter_min_1/in
+ mux_2to1_logic_1/DinB buffer_no_inv_x05
Xbuffer_no_inv_x05_6 avss1p8 mux_2to1_logic_1/DinB avdd1p8 buffer_no_inv_x05_6/inverter_min_1/in
+ buffer_no_inv_x05_7/in buffer_no_inv_x05
Xbuffer_no_inv_x05_7 avss1p8 buffer_no_inv_x05_7/in avdd1p8 buffer_no_inv_x05_7/inverter_min_1/in
+ mux_2to1_logic_3/DinA buffer_no_inv_x05
C0 reg0 mux_2to1_logic_6/sel_b 0.06fF
C1 mux_2to1_logic_4/out mux_2to1_logic_5/out 0.45fF
C2 mux_2to1_logic_2/sel_b mux_2to1_logic_0/out 0.15fF
C3 mux_2to1_logic_6/sel_b mux_2to1_logic_4/DinA 0.01fF
C4 avdd1p8 reg1 0.08fF
C5 mux_2to1_logic_0/DinB mux_2to1_logic_0/sel_b 0.06fF
C6 reg2 mux_2to1_logic_3/DinA 0.33fF
C7 reg2 mux_2to1_logic_1/DinA 0.18fF
C8 buffer_no_inv_x05_13/in clk 0.07fF
C9 mux_2to1_logic_2/out reg0 0.44fF
C10 mux_2to1_logic_4/DinB mux_2to1_logic_3/out 0.18fF
C11 mux_2to1_logic_4/DinB buffer_no_inv_x05_13/inverter_min_1/in 0.11fF
C12 buffer_no_inv_x05_9/in buffer_no_inv_x05_8/inverter_min_1/in 0.07fF
C13 buffer_no_inv_x05_7/in buffer_no_inv_x05_7/inverter_min_1/in 0.12fF
C14 mux_2to1_logic_4/out avdd1p8 0.76fF
C15 mux_2to1_logic_1/DinA mux_2to1_logic_1/out 0.05fF
C16 mux_2to1_logic_4/sel_b mux_2to1_logic_3/DinB 0.04fF
C17 mux_2to1_logic_3/out mux_2to1_logic_3/DinA 0.05fF
C18 mux_2to1_logic_4/DinB reg1 0.40fF
C19 mux_2to1_logic_1/DinB mux_2to1_logic_0/out 0.12fF
C20 buffer_no_inv_x05_11/in buffer_no_inv_x05_10/inverter_min_1/in 0.07fF
C21 avdd1p8 mux_2to1_logic_4/sel_b 0.07fF
C22 mux_2to1_logic_6/sel_b mux_2to1_logic_5/out 0.20fF
C23 buffer_no_inv_x05_3/in mux_2to1_logic_1/DinA 0.16fF
C24 avdd1p8 buffer_no_inv_x05_12/inverter_min_1/in 0.03fF
C25 avdd1p8 buffer_no_inv_x05_11/inverter_min_1/in 0.03fF
C26 reg2 mux_2to1_logic_3/out 0.36fF
C27 mux_2to1_logic_2/out nand_logic_0/in1 0.06fF
C28 reg2 mux_2to1_logic_0/sel_b 0.14fF
C29 mux_2to1_logic_2/sel_b buffer_no_inv_x05_5/in 0.01fF
C30 mux_2to1_logic_4/DinA clk 0.01fF
C31 mux_2to1_logic_3/sel_b mux_2to1_logic_3/DinB 0.21fF
C32 avdd1p8 mux_2to1_logic_0/out 0.43fF
C33 mux_2to1_logic_2/out mux_2to1_logic_5/out 1.29fF
C34 buffer_no_inv_x05_5/in buffer_no_inv_x05_4/inverter_min_1/in 0.07fF
C35 reg2 reg1 2.15fF
C36 mux_2to1_logic_4/out mux_2to1_logic_4/DinB 0.65fF
C37 mux_2to1_logic_3/sel_b avdd1p8 0.09fF
C38 mux_2to1_logic_3/DinB buffer_no_inv_x05_7/inverter_min_1/in 0.10fF
C39 avdd1p8 mux_2to1_logic_6/sel_b 0.05fF
C40 mux_2to1_logic_4/DinB mux_2to1_logic_4/sel_b 0.20fF
C41 mux_2to1_logic_3/DinB mux_2to1_logic_5/sel_b 0.01fF
C42 mux_2to1_logic_4/DinB buffer_no_inv_x05_12/inverter_min_1/in 0.07fF
C43 mux_2to1_logic_0/DinB mux_2to1_logic_0/out 0.14fF
C44 avdd1p8 buffer_no_inv_x05_7/inverter_min_1/in 0.04fF
C45 mux_2to1_logic_1/out reg1 0.36fF
C46 avdd1p8 mux_2to1_logic_5/sel_b 0.09fF
C47 avdd1p8 buffer_no_inv_x05_13/in 0.10fF
C48 buffer_no_inv_x05_9/in mux_2to1_logic_3/DinB 0.10fF
C49 mux_2to1_logic_3/out reg1 0.47fF
C50 mux_2to1_logic_2/out avdd1p8 0.41fF
C51 reg0 mux_2to1_logic_5/out 0.23fF
C52 buffer_no_inv_x05_5/in mux_2to1_logic_1/DinB 0.15fF
C53 mux_2to1_logic_1/DinB mux_2to1_logic_1/sel_b -0.06fF
C54 avdd1p8 buffer_no_inv_x05_9/in 0.10fF
C55 mux_2to1_logic_4/DinA mux_2to1_logic_5/out 0.23fF
C56 mux_2to1_logic_3/sel_b buffer_no_inv_x05_6/inverter_min_1/in 0.01fF
C57 reg2 mux_2to1_logic_4/sel_b 0.06fF
C58 mux_2to1_logic_4/DinB mux_2to1_logic_6/sel_b 0.28fF
C59 mux_2to1_logic_1/DinB clk 0.01fF
C60 clk_out clk 0.33fF
C61 buffer_no_inv_x05_1/inverter_min_1/in buffer_no_inv_x05_1/in 0.12fF
C62 mux_2to1_logic_3/DinB buffer_no_inv_x05_8/inverter_min_1/in 0.10fF
C63 buffer_no_inv_x05_11/in avdd1p8 0.10fF
C64 mux_2to1_logic_1/sel_b avdd1p8 0.09fF
C65 buffer_no_inv_x05_5/in avdd1p8 0.09fF
C66 mux_2to1_logic_1/DinA mux_2to1_logic_0/out 0.12fF
C67 buffer_no_inv_x05_10/inverter_min_1/in mux_2to1_logic_3/DinB 0.12fF
C68 avdd1p8 buffer_no_inv_x05_1/inverter_min_1/in 0.03fF
C69 mux_2to1_logic_4/out mux_2to1_logic_3/out 1.18fF
C70 mux_2to1_logic_3/DinB clk 0.01fF
C71 mux_2to1_logic_4/DinA mux_2to1_logic_3/DinB 0.90fF
C72 mux_2to1_logic_2/sel_b mux_2to1_logic_1/DinB 0.04fF
C73 mux_2to1_logic_4/DinB buffer_no_inv_x05_13/in 0.11fF
C74 mux_2to1_logic_4/DinB mux_2to1_logic_5/sel_b 0.31fF
C75 reg2 mux_2to1_logic_0/out 0.45fF
C76 nand_logic_0/in1 mux_2to1_logic_5/out 0.38fF
C77 avdd1p8 buffer_no_inv_x05_8/inverter_min_1/in 0.03fF
C78 mux_2to1_logic_1/DinB buffer_no_inv_x05_4/inverter_min_1/in 0.15fF
C79 reg0 avdd1p8 0.05fF
C80 avdd1p8 buffer_no_inv_x05_10/inverter_min_1/in 0.03fF
C81 mux_2to1_logic_2/out mux_2to1_logic_4/DinB 0.07fF
C82 avdd1p8 mux_2to1_logic_4/DinA 1.95fF
C83 mux_2to1_logic_4/sel_b mux_2to1_logic_3/out 0.23fF
C84 avdd1p8 clk 1.01fF
C85 mux_2to1_logic_3/sel_b reg2 0.13fF
C86 buffer_no_inv_x05_7/inverter_min_1/in mux_2to1_logic_3/DinA 0.21fF
C87 buffer_no_inv_x05_7/in mux_2to1_logic_3/DinB 0.10fF
C88 mux_2to1_logic_0/DinB mux_2to1_logic_1/sel_b 0.04fF
C89 mux_2to1_logic_0/DinB buffer_no_inv_x05_1/inverter_min_1/in 0.08fF
C90 mux_2to1_logic_4/out reg1 0.37fF
C91 buffer_no_inv_x05_0/inverter_min_1/in buffer_no_inv_x05_1/in 0.07fF
C92 mux_2to1_logic_1/out mux_2to1_logic_0/out 1.27fF
C93 mux_2to1_logic_2/sel_b avdd1p8 0.07fF
C94 avdd1p8 buffer_no_inv_x05_7/in 0.09fF
C95 buffer_no_inv_x05_0/inverter_min_1/in avdd1p8 0.01fF
C96 avdd1p8 buffer_no_inv_x05_4/inverter_min_1/in 0.03fF
C97 mux_2to1_logic_0/DinB clk 0.01fF
C98 mux_2to1_logic_3/sel_b mux_2to1_logic_1/out 0.04fF
C99 mux_2to1_logic_1/DinB buffer_no_inv_x05_3/inverter_min_1/in 0.15fF
C100 buffer_no_inv_x05_5/in buffer_no_inv_x05_5/inverter_min_1/in 0.12fF
C101 mux_2to1_logic_2/out reg2 0.85fF
C102 reg0 mux_2to1_logic_4/DinB -0.24fF
C103 mux_2to1_logic_4/DinB mux_2to1_logic_4/DinA 1.68fF
C104 mux_2to1_logic_4/DinB clk 0.12fF
C105 avdd1p8 buffer_no_inv_x05_2/inverter_min_1/in 0.03fF
C106 buffer_no_inv_x05_9/inverter_min_1/in buffer_no_inv_x05_9/in 0.12fF
C107 avdd1p8 mux_2to1_logic_5/out 0.64fF
C108 reg1 mux_2to1_logic_0/out 0.63fF
C109 mux_2to1_logic_2/out mux_2to1_logic_1/out 0.35fF
C110 avdd1p8 buffer_no_inv_x05_3/inverter_min_1/in 0.03fF
C111 buffer_no_inv_x05_7/in buffer_no_inv_x05_6/inverter_min_1/in 0.07fF
C112 buffer_no_inv_x05_8/inverter_min_1/in mux_2to1_logic_3/DinA 0.12fF
C113 mux_2to1_logic_3/out mux_2to1_logic_5/sel_b 0.37fF
C114 buffer_no_inv_x05_13/inverter_min_1/in buffer_no_inv_x05_13/in 0.12fF
C115 reg2 mux_2to1_logic_1/sel_b 0.13fF
C116 mux_2to1_logic_1/DinB avdd1p8 1.09fF
C117 clk mux_2to1_logic_3/DinA 0.01fF
C118 mux_2to1_logic_4/DinA mux_2to1_logic_3/DinA 0.07fF
C119 mux_2to1_logic_2/out mux_2to1_logic_3/out 0.99fF
C120 avdd1p8 clk_out 0.04fF
C121 mux_2to1_logic_0/DinB buffer_no_inv_x05_2/inverter_min_1/in 0.12fF
C122 mux_2to1_logic_1/DinA clk 0.01fF
C123 reg2 clk 0.12fF
C124 reg2 mux_2to1_logic_4/DinA 0.31fF
C125 avdd1p8 mux_2to1_logic_3/DinB 0.82fF
C126 buffer_no_inv_x05_7/in mux_2to1_logic_3/DinA 0.13fF
C127 avdd1p8 buffer_no_inv_x05_1/in 0.09fF
C128 mux_2to1_logic_5/sel_b reg1 0.06fF
C129 mux_2to1_logic_2/out reg1 1.41fF
C130 mux_2to1_logic_1/DinA buffer_no_inv_x05_4/inverter_min_1/in 0.12fF
C131 mux_2to1_logic_4/DinB mux_2to1_logic_5/out 0.52fF
C132 mux_2to1_logic_2/sel_b reg2 0.07fF
C133 buffer_no_inv_x05_3/in mux_2to1_logic_1/sel_b 0.01fF
C134 mux_2to1_logic_4/out mux_2to1_logic_6/sel_b 0.04fF
C135 mux_2to1_logic_1/DinB buffer_no_inv_x05_6/inverter_min_1/in 0.12fF
C136 buffer_no_inv_x05_1/inverter_min_1/in mux_2to1_logic_0/sel_b 0.01fF
C137 mux_2to1_logic_1/DinB buffer_no_inv_x05_5/inverter_min_1/in 0.23fF
C138 mux_2to1_logic_0/DinB avdd1p8 1.33fF
C139 mux_2to1_logic_4/DinA mux_2to1_logic_3/out 0.12fF
C140 mux_2to1_logic_3/DinB buffer_no_inv_x05_6/inverter_min_1/in 0.02fF
C141 mux_2to1_logic_4/out mux_2to1_logic_5/sel_b 0.20fF
C142 mux_2to1_logic_2/sel_b mux_2to1_logic_1/out 0.19fF
C143 mux_2to1_logic_1/DinA buffer_no_inv_x05_2/inverter_min_1/in 0.10fF
C144 mux_2to1_logic_4/DinB mux_2to1_logic_3/DinB 0.29fF
C145 mux_2to1_logic_4/out mux_2to1_logic_2/out 0.26fF
C146 mux_2to1_logic_1/DinA buffer_no_inv_x05_3/inverter_min_1/in 0.23fF
C147 mux_2to1_logic_1/DinB mux_2to1_logic_3/DinA 0.07fF
C148 avdd1p8 buffer_no_inv_x05_6/inverter_min_1/in 0.03fF
C149 reg0 reg1 0.01fF
C150 mux_2to1_logic_1/DinB mux_2to1_logic_1/DinA 0.66fF
C151 mux_2to1_logic_4/DinB avdd1p8 2.49fF
C152 buffer_no_inv_x05_13/in buffer_no_inv_x05_12/inverter_min_1/in 0.07fF
C153 avdd1p8 buffer_no_inv_x05_5/inverter_min_1/in 0.03fF
C154 mux_2to1_logic_2/out mux_2to1_logic_4/sel_b 0.22fF
C155 reg2 mux_2to1_logic_1/DinB 0.07fF
C156 mux_2to1_logic_3/DinB mux_2to1_logic_3/DinA 1.18fF
C157 mux_2to1_logic_2/sel_b reg1 0.06fF
C158 avdd1p8 mux_2to1_logic_3/DinA 0.81fF
C159 reg2 mux_2to1_logic_3/DinB 0.08fF
C160 buffer_no_inv_x05_4/inverter_min_1/in reg1 0.01fF
C161 reg2 buffer_no_inv_x05_1/in 0.01fF
C162 avdd1p8 mux_2to1_logic_1/DinA 0.55fF
C163 mux_2to1_logic_3/out mux_2to1_logic_5/out 0.07fF
C164 mux_2to1_logic_2/out mux_2to1_logic_0/out 0.05fF
C165 buffer_no_inv_x05_3/in buffer_no_inv_x05_2/inverter_min_1/in 0.07fF
C166 mux_2to1_logic_1/DinB mux_2to1_logic_1/out 0.23fF
C167 reg2 avdd1p8 0.14fF
C168 buffer_no_inv_x05_9/inverter_min_1/in mux_2to1_logic_3/DinB 0.18fF
C169 buffer_no_inv_x05_11/in buffer_no_inv_x05_11/inverter_min_1/in 0.14fF
C170 buffer_no_inv_x05_3/in buffer_no_inv_x05_3/inverter_min_1/in 0.12fF
C171 mux_2to1_logic_4/out mux_2to1_logic_4/DinA 0.27fF
C172 mux_2to1_logic_3/sel_b mux_2to1_logic_2/out 0.33fF
C173 mux_2to1_logic_4/sel_b buffer_no_inv_x05_8/inverter_min_1/in 0.01fF
C174 buffer_no_inv_x05_3/in mux_2to1_logic_1/DinB 0.03fF
C175 buffer_no_inv_x05_9/inverter_min_1/in avdd1p8 0.03fF
C176 mux_2to1_logic_2/out mux_2to1_logic_6/sel_b 0.31fF
C177 mux_2to1_logic_0/DinB mux_2to1_logic_1/DinA 0.11fF
C178 reg0 buffer_no_inv_x05_11/inverter_min_1/in 0.01fF
C179 reg2 mux_2to1_logic_0/DinB 0.06fF
C180 mux_2to1_logic_4/DinA buffer_no_inv_x05_12/inverter_min_1/in 0.12fF
C181 mux_2to1_logic_4/DinA buffer_no_inv_x05_11/inverter_min_1/in 0.08fF
C182 mux_2to1_logic_3/DinB mux_2to1_logic_3/out 0.13fF
C183 avdd1p8 mux_2to1_logic_1/out 0.84fF
C184 buffer_no_inv_x05_6/inverter_min_1/in mux_2to1_logic_3/DinA 0.04fF
C185 nand_logic_0/m1_21_n341# clk_out 0.02fF
C186 mux_2to1_logic_1/sel_b mux_2to1_logic_0/out 0.26fF
C187 mux_2to1_logic_2/out mux_2to1_logic_5/sel_b 0.20fF
C188 avdd1p8 mux_2to1_logic_3/out 0.39fF
C189 buffer_no_inv_x05_13/inverter_min_1/in avdd1p8 0.03fF
C190 buffer_no_inv_x05_3/in avdd1p8 0.11fF
C191 avdd1p8 mux_2to1_logic_0/sel_b 0.05fF
C192 clk mux_2to1_logic_0/out 0.05fF
C193 reg2 mux_2to1_logic_4/DinB 0.05fF
C194 buffer_no_inv_x05_7/in avss1p8 1.12fF
C195 mux_2to1_logic_3/DinA avss1p8 0.02fF
C196 buffer_no_inv_x05_7/inverter_min_1/in avss1p8 1.05fF
C197 buffer_no_inv_x05_6/inverter_min_1/in avss1p8 1.04fF
C198 buffer_no_inv_x05_5/in avss1p8 1.12fF
C199 buffer_no_inv_x05_5/inverter_min_1/in avss1p8 1.04fF
C200 buffer_no_inv_x05_4/inverter_min_1/in avss1p8 1.04fF
C201 buffer_no_inv_x05_3/in avss1p8 1.13fF
C202 buffer_no_inv_x05_3/inverter_min_1/in avss1p8 1.04fF
C203 buffer_no_inv_x05_1/in avss1p8 1.12fF
C204 buffer_no_inv_x05_1/inverter_min_1/in avss1p8 1.04fF
C205 buffer_no_inv_x05_2/inverter_min_1/in avss1p8 1.05fF
C206 clk avss1p8 2.54fF
C207 buffer_no_inv_x05_0/inverter_min_1/in avss1p8 1.03fF
C208 buffer_no_inv_x05_13/in avss1p8 1.12fF
C209 mux_2to1_logic_4/DinB avss1p8 -7.83fF
C210 buffer_no_inv_x05_13/inverter_min_1/in avss1p8 1.04fF
C211 buffer_no_inv_x05_12/inverter_min_1/in avss1p8 1.04fF
C212 buffer_no_inv_x05_11/in avss1p8 1.12fF
C213 buffer_no_inv_x05_11/inverter_min_1/in avss1p8 1.04fF
C214 nand_logic_0/m1_21_n341# avss1p8 0.72fF
C215 clk_out avss1p8 0.27fF
C216 buffer_no_inv_x05_10/inverter_min_1/in avss1p8 1.04fF
C217 nand_logic_0/in1 avss1p8 1.63fF
C218 mux_2to1_logic_6/sel_b avss1p8 2.08fF
C219 reg0 avss1p8 3.16fF
C220 mux_2to1_logic_5/out avss1p8 -1.59fF
C221 mux_2to1_logic_5/sel_b avss1p8 2.05fF
C222 mux_2to1_logic_4/DinA avss1p8 -2.53fF
C223 mux_2to1_logic_4/out avss1p8 -2.14fF
C224 mux_2to1_logic_4/sel_b avss1p8 2.05fF
C225 mux_2to1_logic_3/out avss1p8 -2.13fF
C226 mux_2to1_logic_3/DinB avss1p8 -4.89fF
C227 mux_2to1_logic_3/sel_b avss1p8 2.05fF
C228 mux_2to1_logic_2/out avss1p8 -1.34fF
C229 mux_2to1_logic_2/sel_b avss1p8 2.05fF
C230 reg1 avss1p8 4.95fF
C231 mux_2to1_logic_1/DinA avss1p8 0.68fF
C232 mux_2to1_logic_1/out avss1p8 -2.38fF
C233 mux_2to1_logic_1/DinB avss1p8 -3.84fF
C234 mux_2to1_logic_1/sel_b avss1p8 2.05fF
C235 reg2 avss1p8 13.29fF
C236 avdd1p8 avss1p8 125.49fF
C237 mux_2to1_logic_0/out avss1p8 0.32fF
C238 mux_2to1_logic_0/DinB avss1p8 -0.89fF
C239 mux_2to1_logic_0/sel_b avss1p8 2.04fF
C240 buffer_no_inv_x05_9/in avss1p8 1.12fF
C241 buffer_no_inv_x05_9/inverter_min_1/in avss1p8 1.04fF
C242 buffer_no_inv_x05_8/inverter_min_1/in avss1p8 1.04fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_72JNYZ a_n81_n100# w_n311_n310# a_n128_122# a_111_n100#
+ a_15_n100# a_n173_n100#
X0 a_15_n100# a_n128_122# a_n81_n100# w_n311_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n81_n100# a_n128_122# a_n173_n100# w_n311_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_111_n100# a_n128_122# a_15_n100# w_n311_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_n128_122# a_n81_n100# 0.10fF
C1 a_15_n100# a_111_n100# 0.29fF
C2 a_15_n100# a_n81_n100# 0.29fF
C3 a_n81_n100# a_111_n100# 0.11fF
C4 a_15_n100# a_n173_n100# 0.11fF
C5 a_15_n100# a_n128_122# 0.10fF
C6 a_111_n100# a_n173_n100# 0.06fF
C7 a_n81_n100# a_n173_n100# 0.29fF
C8 a_111_n100# w_n311_n310# 0.15fF
C9 a_15_n100# w_n311_n310# 0.11fF
C10 a_n81_n100# w_n311_n310# 0.11fF
C11 a_n173_n100# w_n311_n310# 0.15fF
C12 a_n128_122# w_n311_n310# 0.49fF
.ends

.subckt sky130_fd_pr__pfet_01v8_2XL9AN VSUBS w_n311_n319# a_n81_n100# a_111_n100#
+ a_n129_131# a_15_n100# a_n173_n100#
X0 a_15_n100# a_n129_131# a_n81_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_n100# a_n129_131# a_15_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n81_n100# a_n129_131# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 w_n311_n319# a_n173_n100# 0.12fF
C1 a_n81_n100# a_15_n100# 0.29fF
C2 a_111_n100# w_n311_n319# 0.12fF
C3 a_n81_n100# a_n173_n100# 0.29fF
C4 w_n311_n319# a_n129_131# 0.16fF
C5 a_n173_n100# a_15_n100# 0.11fF
C6 a_111_n100# a_n81_n100# 0.11fF
C7 a_n81_n100# a_n129_131# 0.08fF
C8 a_n81_n100# w_n311_n319# 0.08fF
C9 a_111_n100# a_15_n100# 0.29fF
C10 a_15_n100# a_n129_131# 0.08fF
C11 w_n311_n319# a_15_n100# 0.08fF
C12 a_111_n100# a_n173_n100# 0.06fF
C13 a_111_n100# VSUBS 0.03fF
C14 a_15_n100# VSUBS 0.03fF
C15 a_n81_n100# VSUBS 0.03fF
C16 a_n173_n100# VSUBS 0.03fF
C17 a_n129_131# VSUBS 0.32fF
C18 w_n311_n319# VSUBS 2.34fF
.ends

.subckt sky130_fd_pr__pfet_01v8_2XUYGK VSUBS a_n269_n100# a_n81_n100# w_n407_n319#
+ a_111_n100# a_n177_n100# a_15_n100# a_207_n100# a_n225_131#
X0 a_207_n100# a_n225_131# a_111_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_15_n100# a_n225_131# a_n81_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_111_n100# a_n225_131# a_15_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n81_n100# a_n225_131# a_n177_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n177_n100# a_n225_131# a_n269_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_111_n100# a_n81_n100# 0.11fF
C1 w_n407_n319# a_n269_n100# 0.10fF
C2 a_n177_n100# a_n81_n100# 0.29fF
C3 a_111_n100# a_n269_n100# 0.05fF
C4 a_15_n100# a_n225_131# 0.08fF
C5 a_15_n100# w_n407_n319# 0.06fF
C6 a_n177_n100# a_n269_n100# 0.29fF
C7 w_n407_n319# a_n225_131# 0.25fF
C8 a_15_n100# a_207_n100# 0.11fF
C9 a_15_n100# a_111_n100# 0.29fF
C10 a_111_n100# a_n225_131# 0.08fF
C11 w_n407_n319# a_207_n100# 0.10fF
C12 a_n269_n100# a_n81_n100# 0.11fF
C13 a_15_n100# a_n177_n100# 0.11fF
C14 w_n407_n319# a_111_n100# 0.05fF
C15 a_n177_n100# a_n225_131# 0.08fF
C16 a_111_n100# a_207_n100# 0.29fF
C17 a_n177_n100# w_n407_n319# 0.05fF
C18 a_n177_n100# a_207_n100# 0.05fF
C19 a_15_n100# a_n81_n100# 0.29fF
C20 a_n81_n100# a_n225_131# 0.08fF
C21 a_n177_n100# a_111_n100# 0.06fF
C22 w_n407_n319# a_n81_n100# 0.06fF
C23 a_15_n100# a_n269_n100# 0.06fF
C24 a_n81_n100# a_207_n100# 0.06fF
C25 a_207_n100# VSUBS 0.03fF
C26 a_111_n100# VSUBS 0.03fF
C27 a_15_n100# VSUBS 0.03fF
C28 a_n81_n100# VSUBS 0.03fF
C29 a_n177_n100# VSUBS 0.03fF
C30 a_n269_n100# VSUBS 0.03fF
C31 a_n225_131# VSUBS 0.54fF
C32 w_n407_n319# VSUBS 2.92fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_2AP43D a_15_n81# a_n33_41# w_n211_n229# a_n73_n81#
X0 a_15_n81# a_n33_41# a_n73_n81# w_n211_n229# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
C0 a_n73_n81# a_n33_41# 0.02fF
C1 a_n33_41# a_15_n81# 0.02fF
C2 a_n73_n81# a_15_n81# 0.17fF
C3 a_15_n81# w_n211_n229# 0.12fF
C4 a_n73_n81# w_n211_n229# 0.12fF
C5 a_n33_41# w_n211_n229# 0.18fF
.ends

.subckt res_amp_lin clk vctrl avdd1p8 avss1p8 a_3747_261# vp inn outn outp inp
Xsky130_fd_pr__pfet_01v8_2XL9AN_0 avss1p8 avdd1p8 a_3747_261# a_3747_261# clk avdd1p8
+ avdd1p8 sky130_fd_pr__pfet_01v8_2XL9AN
Xsky130_fd_pr__pfet_01v8_2XUYGK_0 avss1p8 a_3747_261# a_3747_261# avdd1p8 a_3747_261#
+ vp vp vp vctrl sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_1 avss1p8 vp vp avdd1p8 vp outp outp outp inn sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__nfet_01v8_lvt_2AP43D_0 avss1p8 clk avss1p8 outp sky130_fd_pr__nfet_01v8_lvt_2AP43D
Xsky130_fd_pr__pfet_01v8_2XUYGK_2 avss1p8 vp vp avdd1p8 vp outp outp outp inn sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__nfet_01v8_lvt_2AP43D_1 avss1p8 clk avss1p8 outn sky130_fd_pr__nfet_01v8_lvt_2AP43D
Xsky130_fd_pr__pfet_01v8_2XUYGK_3 avss1p8 vp vp avdd1p8 vp outn outn outn inp sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_4 avss1p8 vp vp avdd1p8 vp outn outn outn inp sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_5 avss1p8 vp vp avdd1p8 vp outp outp outp inn sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_6 avss1p8 vp vp avdd1p8 vp outp outp outp inn sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_7 avss1p8 vp vp avdd1p8 vp outn outn outn inp sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_8 avss1p8 vp vp avdd1p8 vp outn outn outn inp sky130_fd_pr__pfet_01v8_2XUYGK
C0 avdd1p8 outp 1.56fF
C1 clk vctrl 0.02fF
C2 inp outp 1.28fF
C3 outn inn 1.15fF
C4 vp outn 4.23fF
C5 clk outn 0.71fF
C6 avdd1p8 vctrl 1.19fF
C7 avdd1p8 outn 1.33fF
C8 vp inn 0.84fF
C9 clk vp 0.79fF
C10 a_3747_261# vctrl 0.76fF
C11 inp outn 5.59fF
C12 avdd1p8 inn 1.05fF
C13 avdd1p8 vp 6.92fF
C14 avdd1p8 clk 2.36fF
C15 inp inn 2.67fF
C16 vp inp 0.78fF
C17 clk inp 0.06fF
C18 outn outp 4.18fF
C19 vp a_3747_261# 1.08fF
C20 clk a_3747_261# 0.44fF
C21 avdd1p8 inp 1.02fF
C22 avdd1p8 a_3747_261# 1.24fF
C23 inn outp 5.76fF
C24 vp outp 4.81fF
C25 clk outp 0.56fF
C26 outn avss1p8 0.69fF
C27 inp avss1p8 -0.11fF
C28 outp avss1p8 -0.62fF
C29 vp avss1p8 -4.89fF
C30 inn avss1p8 0.23fF
C31 avdd1p8 avss1p8 31.50fF
C32 clk avss1p8 1.49fF
C33 a_3747_261# avss1p8 -0.95fF
C34 vctrl avss1p8 -0.82fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_595QY5 a_n269_n100# a_n81_n100# a_111_n100# a_n177_n100#
+ a_15_n100# w_n407_n310# a_207_n100# a_n225_n188#
X0 a_207_n100# a_n225_n188# a_111_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_15_n100# a_n225_n188# a_n81_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n81_n100# a_n225_n188# a_n177_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_111_n100# a_n225_n188# a_15_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n177_n100# a_n225_n188# a_n269_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_n225_n188# a_n177_n100# 0.10fF
C1 a_n81_n100# a_15_n100# 0.29fF
C2 a_111_n100# a_n177_n100# 0.06fF
C3 a_n269_n100# a_n177_n100# 0.29fF
C4 a_n225_n188# a_15_n100# 0.10fF
C5 a_111_n100# a_15_n100# 0.29fF
C6 a_n269_n100# a_15_n100# 0.06fF
C7 a_n225_n188# a_n81_n100# 0.10fF
C8 a_111_n100# a_n81_n100# 0.11fF
C9 a_207_n100# a_n177_n100# 0.05fF
C10 a_n269_n100# a_n81_n100# 0.11fF
C11 a_n225_n188# a_111_n100# 0.10fF
C12 a_207_n100# a_15_n100# 0.11fF
C13 a_n269_n100# a_111_n100# 0.05fF
C14 a_207_n100# a_n81_n100# 0.06fF
C15 a_n177_n100# a_15_n100# 0.11fF
C16 a_n177_n100# a_n81_n100# 0.29fF
C17 a_207_n100# a_111_n100# 0.29fF
C18 a_207_n100# w_n407_n310# 0.13fF
C19 a_111_n100# w_n407_n310# 0.08fF
C20 a_15_n100# w_n407_n310# 0.09fF
C21 a_n81_n100# w_n407_n310# 0.09fF
C22 a_n177_n100# w_n407_n310# 0.08fF
C23 a_n269_n100# w_n407_n310# 0.13fF
C24 a_n225_n188# w_n407_n310# 0.80fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_9B2JY7 a_n317_n100# a_n33_n100# a_n225_n100# a_n271_122#
+ a_63_n100# a_n129_n100# w_n455_n310# a_255_n100# a_159_n100#
X0 a_63_n100# a_n271_122# a_n33_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n271_122# a_n129_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_159_n100# a_n271_122# a_63_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_255_n100# a_n271_122# a_159_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n225_n100# a_n271_122# a_n317_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n129_n100# a_n271_122# a_n225_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_159_n100# a_63_n100# 0.29fF
C1 a_n317_n100# a_n33_n100# 0.06fF
C2 a_n129_n100# a_n225_n100# 0.29fF
C3 a_159_n100# a_n33_n100# 0.11fF
C4 a_n129_n100# a_63_n100# 0.11fF
C5 a_n225_n100# a_63_n100# 0.06fF
C6 a_n129_n100# a_n33_n100# 0.29fF
C7 a_n271_122# a_159_n100# 0.10fF
C8 a_n225_n100# a_n33_n100# 0.11fF
C9 a_159_n100# a_255_n100# 0.29fF
C10 a_n33_n100# a_63_n100# 0.29fF
C11 a_n271_122# a_n129_n100# 0.10fF
C12 a_n129_n100# a_255_n100# 0.05fF
C13 a_n271_122# a_n225_n100# 0.10fF
C14 a_n271_122# a_63_n100# 0.10fF
C15 a_255_n100# a_63_n100# 0.11fF
C16 a_n317_n100# a_n129_n100# 0.11fF
C17 a_159_n100# a_n129_n100# 0.06fF
C18 a_n317_n100# a_n225_n100# 0.29fF
C19 a_n271_122# a_n33_n100# 0.10fF
C20 a_n33_n100# a_255_n100# 0.06fF
C21 a_159_n100# a_n225_n100# 0.05fF
C22 a_n317_n100# a_63_n100# 0.05fF
C23 a_255_n100# w_n455_n310# 0.13fF
C24 a_159_n100# w_n455_n310# 0.08fF
C25 a_63_n100# w_n455_n310# 0.07fF
C26 a_n33_n100# w_n455_n310# 0.08fF
C27 a_n129_n100# w_n455_n310# 0.07fF
C28 a_n225_n100# w_n455_n310# 0.08fF
C29 a_n317_n100# w_n455_n310# 0.13fF
C30 a_n271_122# w_n455_n310# 0.95fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_MVT43V a_n33_n100# w_n263_n310# a_63_n100# a_n79_122#
+ a_n125_n100#
X0 a_63_n100# a_n79_122# a_n33_n100# w_n263_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n79_122# a_n125_n100# w_n263_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_63_n100# a_n33_n100# 0.29fF
C1 a_n79_122# a_n33_n100# 0.11fF
C2 a_63_n100# a_n125_n100# 0.11fF
C3 a_n79_122# a_n125_n100# 0.02fF
C4 a_n125_n100# a_n33_n100# 0.29fF
C5 a_n79_122# a_63_n100# 0.02fF
C6 a_63_n100# w_n263_n310# 0.16fF
C7 a_n33_n100# w_n263_n310# 0.12fF
C8 a_n125_n100# w_n263_n310# 0.16fF
C9 a_n79_122# w_n263_n310# 0.37fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_NMSMYT a_n33_n100# a_n321_n100# a_n225_n100# w_n551_n310#
+ a_63_n100# a_n368_122# a_n129_n100# a_351_n100# a_255_n100# a_n413_n100# a_159_n100#
X0 a_63_n100# a_n368_122# a_n33_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n368_122# a_n129_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_159_n100# a_n368_122# a_63_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_255_n100# a_n368_122# a_159_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_351_n100# a_n368_122# a_255_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n321_n100# a_n368_122# a_n413_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n225_n100# a_n368_122# a_n321_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n129_n100# a_n368_122# a_n225_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_n225_n100# a_n321_n100# 0.29fF
C1 a_n368_122# a_n33_n100# 0.10fF
C2 a_159_n100# a_255_n100# 0.29fF
C3 a_n321_n100# a_n33_n100# 0.06fF
C4 a_n368_122# a_n321_n100# 0.10fF
C5 a_63_n100# a_n129_n100# 0.11fF
C6 a_n225_n100# a_n129_n100# 0.29fF
C7 a_351_n100# a_255_n100# 0.29fF
C8 a_159_n100# a_351_n100# 0.11fF
C9 a_n33_n100# a_n129_n100# 0.29fF
C10 a_63_n100# a_255_n100# 0.11fF
C11 a_159_n100# a_63_n100# 0.29fF
C12 a_n225_n100# a_n413_n100# 0.11fF
C13 a_n368_122# a_n129_n100# 0.10fF
C14 a_159_n100# a_n225_n100# 0.05fF
C15 a_n413_n100# a_n33_n100# 0.05fF
C16 a_n33_n100# a_255_n100# 0.06fF
C17 a_n321_n100# a_n129_n100# 0.11fF
C18 a_159_n100# a_n33_n100# 0.11fF
C19 a_351_n100# a_63_n100# 0.06fF
C20 a_n368_122# a_255_n100# 0.10fF
C21 a_n368_122# a_159_n100# 0.10fF
C22 a_n413_n100# a_n321_n100# 0.29fF
C23 a_351_n100# a_n33_n100# 0.05fF
C24 a_n225_n100# a_63_n100# 0.06fF
C25 a_63_n100# a_n33_n100# 0.29fF
C26 a_n225_n100# a_n33_n100# 0.11fF
C27 a_n413_n100# a_n129_n100# 0.06fF
C28 a_n368_122# a_63_n100# 0.10fF
C29 a_255_n100# a_n129_n100# 0.05fF
C30 a_159_n100# a_n129_n100# 0.06fF
C31 a_n368_122# a_n225_n100# 0.10fF
C32 a_63_n100# a_n321_n100# 0.05fF
C33 a_351_n100# w_n551_n310# 0.13fF
C34 a_255_n100# w_n551_n310# 0.08fF
C35 a_159_n100# w_n551_n310# 0.07fF
C36 a_63_n100# w_n551_n310# 0.06fF
C37 a_n33_n100# w_n551_n310# 0.04fF
C38 a_n129_n100# w_n551_n310# 0.06fF
C39 a_n225_n100# w_n551_n310# 0.07fF
C40 a_n321_n100# w_n551_n310# 0.08fF
C41 a_n413_n100# w_n551_n310# 0.13fF
C42 a_n368_122# w_n551_n310# 1.26fF
.ends

.subckt sky130_fd_pr__pfet_01v8_XAYTAL VSUBS w_n311_n319# a_n81_n100# a_n129_n197#
+ a_111_n100# a_15_n100# a_n173_n100#
X0 a_15_n100# a_n129_n197# a_n81_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_n100# a_n129_n197# a_15_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n81_n100# a_n129_n197# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_111_n100# w_n311_n319# 0.12fF
C1 w_n311_n319# a_n173_n100# 0.12fF
C2 a_n81_n100# a_15_n100# 0.29fF
C3 a_111_n100# a_n173_n100# 0.06fF
C4 a_n129_n197# w_n311_n319# 0.17fF
C5 a_n81_n100# w_n311_n319# 0.08fF
C6 a_111_n100# a_n81_n100# 0.11fF
C7 a_n81_n100# a_n173_n100# 0.29fF
C8 a_n81_n100# a_n129_n197# 0.08fF
C9 a_15_n100# w_n311_n319# 0.08fF
C10 a_111_n100# a_15_n100# 0.29fF
C11 a_15_n100# a_n173_n100# 0.11fF
C12 a_n129_n197# a_15_n100# 0.08fF
C13 a_111_n100# VSUBS 0.03fF
C14 a_15_n100# VSUBS 0.03fF
C15 a_n81_n100# VSUBS 0.03fF
C16 a_n173_n100# VSUBS 0.03fF
C17 a_n129_n197# VSUBS 0.34fF
C18 w_n311_n319# VSUBS 2.34fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_B2JNY3 a_n33_n100# a_63_n100# a_n221_n100# a_n129_n100#
+ w_n359_n310# a_n176_122# a_159_n100#
X0 a_63_n100# a_n176_122# a_n33_n100# w_n359_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n176_122# a_n129_n100# w_n359_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_159_n100# a_n176_122# a_63_n100# w_n359_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n129_n100# a_n176_122# a_n221_n100# w_n359_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_n176_122# a_n129_n100# 0.10fF
C1 a_n33_n100# a_63_n100# 0.29fF
C2 a_159_n100# a_n129_n100# 0.06fF
C3 a_159_n100# a_n221_n100# 0.05fF
C4 a_n221_n100# a_n129_n100# 0.29fF
C5 a_n33_n100# a_n176_122# 0.10fF
C6 a_159_n100# a_n33_n100# 0.11fF
C7 a_n33_n100# a_n129_n100# 0.29fF
C8 a_n33_n100# a_n221_n100# 0.11fF
C9 a_63_n100# a_n176_122# 0.10fF
C10 a_159_n100# a_63_n100# 0.29fF
C11 a_63_n100# a_n129_n100# 0.11fF
C12 a_n221_n100# a_63_n100# 0.06fF
C13 a_159_n100# w_n359_n310# 0.13fF
C14 a_63_n100# w_n359_n310# 0.10fF
C15 a_n33_n100# w_n359_n310# 0.10fF
C16 a_n129_n100# w_n359_n310# 0.10fF
C17 a_n221_n100# w_n359_n310# 0.13fF
C18 a_n176_122# w_n359_n310# 0.64fF
.ends

.subckt sky130_fd_pr__pfet_01v8_XACJHL VSUBS a_n81_n197# w_n263_n319# a_n33_n100#
+ a_63_n100# a_n125_n100#
X0 a_63_n100# a_n81_n197# a_n33_n100# w_n263_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n197# a_n125_n100# w_n263_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 w_n263_n319# a_n125_n100# 0.13fF
C1 a_n33_n100# a_63_n100# 0.29fF
C2 a_n81_n197# w_n263_n319# 0.11fF
C3 a_n33_n100# w_n263_n319# 0.09fF
C4 a_n33_n100# a_n125_n100# 0.29fF
C5 a_n33_n100# a_n81_n197# 0.08fF
C6 a_63_n100# w_n263_n319# 0.13fF
C7 a_63_n100# a_n125_n100# 0.11fF
C8 a_63_n100# VSUBS 0.03fF
C9 a_n33_n100# VSUBS 0.03fF
C10 a_n125_n100# VSUBS 0.03fF
C11 a_n81_n197# VSUBS 0.23fF
C12 w_n263_n319# VSUBS 2.05fF
.ends

.subckt iref_ctrl_res_amp m1_n356_n363# avss1p8 vctrl reg2 avdd1p8 reg0 m1_1996_n363#
+ reg1 iref m1_511_801# m1_964_n363# m1_1384_n363#
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_0 iref m1_n356_n363# m1_n356_n363# iref iref iref
+ avss1p8 iref m1_n356_n363# sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_1 avss1p8 m1_n356_n363# m1_n356_n363# avdd1p8
+ avss1p8 avss1p8 avss1p8 avss1p8 m1_n356_n363# sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_MVT43V_0 m1_964_n363# avss1p8 vctrl iref vctrl sky130_fd_pr__nfet_01v8_lvt_MVT43V
Xsky130_fd_pr__nfet_01v8_lvt_MVT43V_1 m1_964_n363# avss1p8 avss1p8 reg0 avss1p8 sky130_fd_pr__nfet_01v8_lvt_MVT43V
Xsky130_fd_pr__nfet_01v8_lvt_NMSMYT_0 vctrl m1_1996_n363# vctrl avss1p8 m1_1996_n363#
+ iref m1_1996_n363# vctrl m1_1996_n363# vctrl vctrl sky130_fd_pr__nfet_01v8_lvt_NMSMYT
Xsky130_fd_pr__nfet_01v8_lvt_NMSMYT_1 avss1p8 m1_1996_n363# avss1p8 avss1p8 m1_1996_n363#
+ reg2 m1_1996_n363# avss1p8 m1_1996_n363# avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt_NMSMYT
Xsky130_fd_pr__nfet_01v8_lvt_72JNYZ_0 m1_448_n363# avss1p8 iref m1_448_n363# vctrl
+ vctrl sky130_fd_pr__nfet_01v8_lvt_72JNYZ
Xsky130_fd_pr__nfet_01v8_lvt_72JNYZ_1 m1_448_n363# avss1p8 avdd1p8 m1_448_n363# avss1p8
+ avss1p8 sky130_fd_pr__nfet_01v8_lvt_72JNYZ
Xsky130_fd_pr__pfet_01v8_XAYTAL_0 avss1p8 avdd1p8 m1_511_801# avss1p8 m1_511_801#
+ avdd1p8 avdd1p8 sky130_fd_pr__pfet_01v8_XAYTAL
Xsky130_fd_pr__nfet_01v8_lvt_B2JNY3_0 vctrl m1_1384_n363# vctrl m1_1384_n363# avss1p8
+ iref vctrl sky130_fd_pr__nfet_01v8_lvt_B2JNY3
Xsky130_fd_pr__nfet_01v8_lvt_B2JNY3_1 avss1p8 m1_1384_n363# avss1p8 m1_1384_n363#
+ avss1p8 reg1 avss1p8 sky130_fd_pr__nfet_01v8_lvt_B2JNY3
Xsky130_fd_pr__pfet_01v8_XACJHL_0 avss1p8 vctrl avdd1p8 m1_511_801# vctrl vctrl sky130_fd_pr__pfet_01v8_XACJHL
C0 m1_1996_n363# reg2 1.30fF
C1 m1_1384_n363# reg1 0.85fF
C2 m1_448_n363# m1_n356_n363# 0.17fF
C3 m1_964_n363# iref 0.11fF
C4 vctrl reg1 0.06fF
C5 m1_964_n363# reg0 0.47fF
C6 iref reg0 0.02fF
C7 iref m1_n356_n363# 1.89fF
C8 m1_448_n363# vctrl 1.16fF
C9 m1_1996_n363# reg1 0.06fF
C10 m1_964_n363# m1_1384_n363# 0.18fF
C11 m1_1384_n363# iref 0.22fF
C12 reg2 reg1 0.04fF
C13 m1_448_n363# avdd1p8 0.77fF
C14 m1_964_n363# vctrl 0.52fF
C15 m1_1384_n363# reg0 0.06fF
C16 vctrl iref 2.27fF
C17 avdd1p8 iref 0.32fF
C18 vctrl reg0 0.04fF
C19 vctrl m1_n356_n363# 0.08fF
C20 m1_511_801# iref 0.05fF
C21 avdd1p8 reg0 0.03fF
C22 avdd1p8 m1_n356_n363# 1.41fF
C23 m1_1996_n363# iref 0.41fF
C24 reg2 iref 0.03fF
C25 m1_1384_n363# vctrl 0.95fF
C26 avdd1p8 vctrl 0.52fF
C27 m1_1996_n363# m1_1384_n363# 0.18fF
C28 m1_511_801# vctrl 1.08fF
C29 avdd1p8 m1_511_801# 1.05fF
C30 m1_1996_n363# vctrl 1.72fF
C31 reg1 iref 0.03fF
C32 vctrl reg2 0.07fF
C33 reg1 reg0 0.04fF
C34 m1_448_n363# m1_964_n363# 0.24fF
C35 m1_448_n363# iref 0.29fF
C36 m1_511_801# avss1p8 -1.62fF
C37 m1_1384_n363# avss1p8 1.30fF
C38 reg1 avss1p8 1.36fF
C39 m1_448_n363# avss1p8 -0.27fF
C40 vctrl avss1p8 2.17fF
C41 m1_1996_n363# avss1p8 -0.61fF
C42 reg2 avss1p8 1.98fF
C43 reg0 avss1p8 0.44fF
C44 m1_964_n363# avss1p8 -0.38fF
C45 avdd1p8 avss1p8 6.02fF
C46 m1_n356_n363# avss1p8 1.89fF
C47 iref avss1p8 2.30fF
.ends

.subckt res_amp_lin_prog delay_cell_buff_0/mux_2to1_logic_0/out iref_ctrl_res_amp_0/m1_964_n363#
+ delay_reg2 avdd1p8 inp delay_cell_buff_0/mux_2to1_logic_3/DinA res_amp_lin_0/vctrl
+ delay_cell_buff_0/mux_2to1_logic_3/out iref_ctrl_res_amp_0/m1_511_801# res_amp_lin_0/clk
+ delay_cell_buff_0/nand_logic_0/in1 outp_cap avss1p8 outn_cap clk delay_cell_buff_0/mux_2to1_logic_1/sel_b
+ delay_reg0 delay_cell_buff_0/mux_2to1_logic_4/DinA delay_cell_buff_0/mux_2to1_logic_4/DinB
+ outn delay_cell_buff_0/mux_2to1_logic_1/DinA outp delay_cell_buff_0/mux_2to1_logic_5/out
+ delay_cell_buff_0/buffer_no_inv_x05_2/inverter_min_1/in delay_cell_buff_0/mux_2to1_logic_3/DinB
+ iref_reg0 delay_cell_buff_0/buffer_no_inv_x05_13/inverter_min_1/in iref_reg1 iref_reg2
+ iref_ctrl_res_amp_0/m1_1384_n363# delay_cell_buff_0/buffer_no_inv_x05_3/in res_amp_lin_0/vp
+ delay_cell_buff_0/nand_logic_0/m1_21_n341# delay_cell_buff_0/mux_2to1_logic_1/out
+ delay_cell_buff_0/mux_2to1_logic_2/out delay_cell_buff_0/buffer_no_inv_x05_12/inverter_min_1/in
+ iref delay_cell_buff_0/buffer_no_inv_x05_7/inverter_min_1/in iref_ctrl_res_amp_0/m1_n356_n363#
+ res_amp_lin_0/a_3747_261# delay_reg1 delay_cell_buff_0/buffer_no_inv_x05_13/in inn
+ delay_cell_buff_0/mux_2to1_logic_4/out iref_ctrl_res_amp_0/m1_1996_n363# delay_cell_buff_0/buffer_no_inv_x05_10/inverter_min_1/in
+ inverter_min_x4_0/out delay_cell_buff_0/mux_2to1_logic_4/sel_b rst
Xsky130_fd_pr__pfet_01v8_lvt_4L9VGG_0 avss1p8 outn_cap avdd1p8 outn_cap res_amp_lin_0/clk
+ outn outn outn outn_cap sky130_fd_pr__pfet_01v8_lvt_4L9VGG
Xsky130_fd_pr__pfet_01v8_lvt_4L9VGG_1 avss1p8 outp_cap avdd1p8 outp_cap res_amp_lin_0/clk
+ outp outp outp outp_cap sky130_fd_pr__pfet_01v8_lvt_4L9VGG
Xdelay_cell_buff_0 delay_cell_buff_0/buffer_no_inv_x05_2/inverter_min_1/in delay_reg2
+ avss1p8 delay_cell_buff_0/mux_2to1_logic_4/DinA avdd1p8 delay_cell_buff_0/buffer_no_inv_x05_13/in
+ clk delay_cell_buff_0/mux_2to1_logic_3/DinA res_amp_lin_0/clk delay_cell_buff_0/mux_2to1_logic_3/DinB
+ delay_reg0 delay_cell_buff_0/buffer_no_inv_x05_10/inverter_min_1/in delay_reg1 delay_cell_buff_0/buffer_no_inv_x05_7/inverter_min_1/in
+ delay_cell_buff_0/nand_logic_0/in1 delay_cell_buff_0/mux_2to1_logic_2/out delay_cell_buff_0/mux_2to1_logic_4/sel_b
+ delay_cell_buff_0/mux_2to1_logic_4/out delay_cell_buff_0/mux_2to1_logic_1/DinA delay_cell_buff_0/mux_2to1_logic_1/sel_b
+ delay_cell_buff_0/buffer_no_inv_x05_3/in delay_cell_buff_0/mux_2to1_logic_5/out
+ delay_cell_buff_0/mux_2to1_logic_0/out delay_cell_buff_0/mux_2to1_logic_4/DinB delay_cell_buff_0/mux_2to1_logic_3/out
+ delay_cell_buff_0/buffer_no_inv_x05_13/inverter_min_1/in delay_cell_buff_0/mux_2to1_logic_1/out
+ avss1p8 delay_cell_buff_0/buffer_no_inv_x05_12/inverter_min_1/in delay_cell_buff_0/nand_logic_0/m1_21_n341#
+ delay_cell_buff
Xinverter_min_x4_0 avdd1p8 res_amp_lin_0/clk avss1p8 inverter_min_x4_0/out inverter_min_x4
Xsky130_fd_pr__nfet_01v8_lvt_72JNYZ_0 outn_cap avss1p8 rst outn_cap avss1p8 avss1p8
+ sky130_fd_pr__nfet_01v8_lvt_72JNYZ
Xres_amp_lin_0 res_amp_lin_0/clk res_amp_lin_0/vctrl avdd1p8 avss1p8 res_amp_lin_0/a_3747_261#
+ res_amp_lin_0/vp inn outn outp inp res_amp_lin
Xsky130_fd_pr__nfet_01v8_lvt_72JNYZ_1 outp_cap avss1p8 rst outp_cap avss1p8 avss1p8
+ sky130_fd_pr__nfet_01v8_lvt_72JNYZ
Xsky130_fd_pr__nfet_01v8_lvt_595QY5_0 outn outn outn outn_cap outn_cap avss1p8 outn_cap
+ inverter_min_x4_0/out sky130_fd_pr__nfet_01v8_lvt_595QY5
Xsky130_fd_pr__nfet_01v8_lvt_595QY5_1 outp outp outp outp_cap outp_cap avss1p8 outp_cap
+ inverter_min_x4_0/out sky130_fd_pr__nfet_01v8_lvt_595QY5
Xiref_ctrl_res_amp_0 iref_ctrl_res_amp_0/m1_n356_n363# avss1p8 res_amp_lin_0/vctrl
+ iref_reg2 avdd1p8 iref_reg0 iref_ctrl_res_amp_0/m1_1996_n363# iref_reg1 iref iref_ctrl_res_amp_0/m1_511_801#
+ iref_ctrl_res_amp_0/m1_964_n363# iref_ctrl_res_amp_0/m1_1384_n363# iref_ctrl_res_amp
C0 outp res_amp_lin_0/clk 0.09fF
C1 inverter_min_x4_0/out rst 0.01fF
C2 avdd1p8 outn_cap 0.26fF
C3 outp_cap avdd1p8 0.25fF
C4 inverter_min_x4_0/out outn_cap 0.57fF
C5 outp_cap inverter_min_x4_0/out 0.57fF
C6 rst outn_cap 0.34fF
C7 outp_cap rst 0.34fF
C8 res_amp_lin_0/clk avdd1p8 1.99fF
C9 avdd1p8 outn 0.36fF
C10 res_amp_lin_0/clk inverter_min_x4_0/out 0.14fF
C11 inverter_min_x4_0/out outn 0.32fF
C12 outp avdd1p8 0.34fF
C13 outp inverter_min_x4_0/out 0.32fF
C14 res_amp_lin_0/clk outn_cap 1.04fF
C15 outn_cap outn 1.90fF
C16 outp_cap res_amp_lin_0/clk 1.04fF
C17 res_amp_lin_0/vctrl iref 0.10fF
C18 res_amp_lin_0/clk outn 0.09fF
C19 avdd1p8 res_amp_lin_0/vctrl 1.42fF
C20 outp_cap outp 1.90fF
C21 iref_ctrl_res_amp_0/m1_511_801# avss1p8 -1.87fF
C22 iref_ctrl_res_amp_0/m1_1384_n363# avss1p8 0.47fF
C23 iref_reg1 avss1p8 0.47fF
C24 iref_ctrl_res_amp_0/m1_448_n363# avss1p8 -1.10fF
C25 res_amp_lin_0/vctrl avss1p8 -1.88fF
C26 iref_ctrl_res_amp_0/m1_1996_n363# avss1p8 -2.23fF
C27 iref_reg2 avss1p8 -0.15fF
C28 iref_reg0 avss1p8 -0.42fF
C29 iref_ctrl_res_amp_0/m1_964_n363# avss1p8 -1.03fF
C30 iref_ctrl_res_amp_0/m1_n356_n363# avss1p8 0.51fF
C31 iref avss1p8 0.07fF
C32 outn avss1p8 1.87fF
C33 inp avss1p8 -0.35fF
C34 outp avss1p8 -4.58fF
C35 res_amp_lin_0/vp avss1p8 -4.89fF
C36 inn avss1p8 0.17fF
C37 res_amp_lin_0/a_3747_261# avss1p8 -0.95fF
C38 outn_cap avss1p8 -1.33fF
C39 rst avss1p8 0.58fF
C40 inverter_min_x4_0/out avss1p8 7.53fF
C41 res_amp_lin_0/clk avss1p8 5.34fF
C42 delay_cell_buff_0/buffer_no_inv_x05_7/in avss1p8 1.07fF
C43 delay_cell_buff_0/mux_2to1_logic_3/DinA avss1p8 -0.04fF
C44 delay_cell_buff_0/buffer_no_inv_x05_7/inverter_min_1/in avss1p8 1.03fF
C45 delay_cell_buff_0/buffer_no_inv_x05_6/inverter_min_1/in avss1p8 1.03fF
C46 delay_cell_buff_0/buffer_no_inv_x05_5/in avss1p8 1.07fF
C47 delay_cell_buff_0/buffer_no_inv_x05_5/inverter_min_1/in avss1p8 1.03fF
C48 delay_cell_buff_0/buffer_no_inv_x05_4/inverter_min_1/in avss1p8 1.03fF
C49 delay_cell_buff_0/buffer_no_inv_x05_3/in avss1p8 1.07fF
C50 delay_cell_buff_0/buffer_no_inv_x05_3/inverter_min_1/in avss1p8 1.03fF
C51 delay_cell_buff_0/buffer_no_inv_x05_1/in avss1p8 1.07fF
C52 delay_cell_buff_0/buffer_no_inv_x05_1/inverter_min_1/in avss1p8 1.03fF
C53 delay_cell_buff_0/buffer_no_inv_x05_2/inverter_min_1/in avss1p8 1.03fF
C54 clk avss1p8 -4.09fF
C55 delay_cell_buff_0/buffer_no_inv_x05_0/inverter_min_1/in avss1p8 1.03fF
C56 delay_cell_buff_0/buffer_no_inv_x05_13/in avss1p8 1.07fF
C57 delay_cell_buff_0/mux_2to1_logic_4/DinB avss1p8 -7.88fF
C58 delay_cell_buff_0/buffer_no_inv_x05_13/inverter_min_1/in avss1p8 1.03fF
C59 delay_cell_buff_0/buffer_no_inv_x05_12/inverter_min_1/in avss1p8 1.03fF
C60 delay_cell_buff_0/buffer_no_inv_x05_11/in avss1p8 1.07fF
C61 delay_cell_buff_0/buffer_no_inv_x05_11/inverter_min_1/in avss1p8 1.03fF
C62 delay_cell_buff_0/nand_logic_0/m1_21_n341# avss1p8 0.72fF
C63 delay_cell_buff_0/buffer_no_inv_x05_10/inverter_min_1/in avss1p8 1.03fF
C64 delay_cell_buff_0/nand_logic_0/in1 avss1p8 1.54fF
C65 delay_cell_buff_0/mux_2to1_logic_6/sel_b avss1p8 2.03fF
C66 delay_reg0 avss1p8 2.77fF
C67 delay_cell_buff_0/mux_2to1_logic_5/out avss1p8 -1.67fF
C68 delay_cell_buff_0/mux_2to1_logic_5/sel_b avss1p8 2.03fF
C69 delay_cell_buff_0/mux_2to1_logic_4/DinA avss1p8 -2.58fF
C70 delay_cell_buff_0/mux_2to1_logic_4/out avss1p8 -2.25fF
C71 delay_cell_buff_0/mux_2to1_logic_4/sel_b avss1p8 2.03fF
C72 delay_cell_buff_0/mux_2to1_logic_3/out avss1p8 -2.69fF
C73 delay_cell_buff_0/mux_2to1_logic_3/DinB avss1p8 -4.96fF
C74 delay_cell_buff_0/mux_2to1_logic_3/sel_b avss1p8 2.03fF
C75 delay_cell_buff_0/mux_2to1_logic_2/out avss1p8 -4.71fF
C76 delay_cell_buff_0/mux_2to1_logic_2/sel_b avss1p8 2.03fF
C77 delay_reg1 avss1p8 3.80fF
C78 delay_cell_buff_0/mux_2to1_logic_1/DinA avss1p8 0.63fF
C79 delay_cell_buff_0/mux_2to1_logic_1/out avss1p8 -2.49fF
C80 delay_cell_buff_0/mux_2to1_logic_1/DinB avss1p8 -3.92fF
C81 delay_cell_buff_0/mux_2to1_logic_1/sel_b avss1p8 2.03fF
C82 delay_reg2 avss1p8 11.07fF
C83 avdd1p8 avss1p8 177.60fF
C84 delay_cell_buff_0/mux_2to1_logic_0/out avss1p8 -0.27fF
C85 delay_cell_buff_0/mux_2to1_logic_0/DinB avss1p8 -0.97fF
C86 delay_cell_buff_0/mux_2to1_logic_0/sel_b avss1p8 2.03fF
C87 delay_cell_buff_0/buffer_no_inv_x05_9/in avss1p8 1.07fF
C88 delay_cell_buff_0/buffer_no_inv_x05_9/inverter_min_1/in avss1p8 1.03fF
C89 delay_cell_buff_0/buffer_no_inv_x05_8/inverter_min_1/in avss1p8 1.03fF
C90 outp_cap avss1p8 -6.93fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_U5ZKVF VSUBS m3_n700_n850# c1_n600_n750#
X0 c1_n600_n750# m3_n700_n850# sky130_fd_pr__cap_mim_m3_1 l=7.5e+06u w=5.5e+06u
C0 c1_n600_n750# m3_n700_n850# 5.48fF
C1 m3_n700_n850# VSUBS 1.98fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_D3F744 VSUBS a_n285_n236# a_355_n236# a_n29_n236#
+ a_n413_n236# a_99_n236# a_n611_n262# a_483_n236# a_n669_n236# w_n807_n384# a_n157_n236#
+ a_n541_n236# a_227_n236# a_611_n236#
X0 a_n157_n236# a_n611_n262# a_n285_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X1 a_611_n236# a_n611_n262# a_483_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X2 a_227_n236# a_n611_n262# a_99_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X3 a_n285_n236# a_n611_n262# a_n413_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X4 a_99_n236# a_n611_n262# a_n29_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X5 a_355_n236# a_n611_n262# a_227_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X6 a_483_n236# a_n611_n262# a_355_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X7 a_n29_n236# a_n611_n262# a_n157_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X8 a_n413_n236# a_n611_n262# a_n541_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X9 a_n541_n236# a_n611_n262# a_n669_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
C0 a_483_n236# a_227_n236# 0.15fF
C1 a_n541_n236# a_n285_n236# 0.15fF
C2 a_n157_n236# a_n541_n236# 0.09fF
C3 a_n413_n236# a_n285_n236# 0.36fF
C4 a_n157_n236# a_n413_n236# 0.15fF
C5 a_n29_n236# a_355_n236# 0.09fF
C6 a_n29_n236# w_n807_n384# 0.02fF
C7 a_355_n236# a_99_n236# 0.15fF
C8 a_n29_n236# a_227_n236# 0.15fF
C9 w_n807_n384# a_99_n236# 0.02fF
C10 a_355_n236# a_611_n236# 0.15fF
C11 a_227_n236# a_99_n236# 0.36fF
C12 w_n807_n384# a_611_n236# 0.19fF
C13 a_n541_n236# a_n413_n236# 0.36fF
C14 a_227_n236# a_611_n236# 0.09fF
C15 a_n669_n236# w_n807_n384# 0.19fF
C16 a_n611_n262# a_355_n236# 0.08fF
C17 a_n611_n262# w_n807_n384# 0.60fF
C18 a_n611_n262# a_227_n236# 0.08fF
C19 a_n29_n236# a_n285_n236# 0.15fF
C20 a_99_n236# a_n285_n236# 0.09fF
C21 a_n29_n236# a_n157_n236# 0.36fF
C22 a_n157_n236# a_99_n236# 0.15fF
C23 a_n669_n236# a_n285_n236# 0.09fF
C24 a_n611_n262# a_n285_n236# 0.08fF
C25 a_355_n236# w_n807_n384# 0.06fF
C26 a_n611_n262# a_n157_n236# 0.08fF
C27 a_355_n236# a_227_n236# 0.36fF
C28 a_227_n236# w_n807_n384# 0.02fF
C29 a_n29_n236# a_n413_n236# 0.09fF
C30 a_n669_n236# a_n541_n236# 0.36fF
C31 a_n611_n262# a_n541_n236# 0.08fF
C32 a_483_n236# a_99_n236# 0.09fF
C33 a_n669_n236# a_n413_n236# 0.15fF
C34 w_n807_n384# a_n285_n236# 0.02fF
C35 a_483_n236# a_611_n236# 0.36fF
C36 a_n611_n262# a_n413_n236# 0.08fF
C37 a_n157_n236# w_n807_n384# 0.02fF
C38 a_n157_n236# a_227_n236# 0.09fF
C39 a_483_n236# a_n611_n262# 0.08fF
C40 a_n29_n236# a_99_n236# 0.36fF
C41 a_n541_n236# w_n807_n384# 0.09fF
C42 a_n157_n236# a_n285_n236# 0.36fF
C43 w_n807_n384# a_n413_n236# 0.06fF
C44 a_n29_n236# a_n611_n262# 0.08fF
C45 a_483_n236# a_355_n236# 0.36fF
C46 a_n611_n262# a_99_n236# 0.08fF
C47 a_483_n236# w_n807_n384# 0.09fF
C48 a_611_n236# VSUBS 0.03fF
C49 a_483_n236# VSUBS 0.03fF
C50 a_355_n236# VSUBS 0.03fF
C51 a_227_n236# VSUBS 0.03fF
C52 a_99_n236# VSUBS 0.03fF
C53 a_n29_n236# VSUBS 0.03fF
C54 a_n157_n236# VSUBS 0.03fF
C55 a_n285_n236# VSUBS 0.03fF
C56 a_n413_n236# VSUBS 0.03fF
C57 a_n541_n236# VSUBS 0.03fF
C58 a_n669_n236# VSUBS 0.03fF
C59 a_n611_n262# VSUBS 1.37fF
C60 w_n807_n384# VSUBS 6.11fF
.ends

.subckt sky130_fd_pr__pfet_01v8_VCU74W VSUBS a_495_n100# a_n81_n100# a_399_n100# a_687_n100#
+ a_n749_n100# a_n273_n100# a_111_n100# a_n177_n100# a_n561_n100# a_15_n100# a_n465_n100#
+ a_n705_n197# a_303_n100# a_n369_n100# w_n887_n319# a_207_n100# a_n657_n100# a_591_n100#
X0 a_303_n100# a_n705_n197# a_207_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_591_n100# a_n705_n197# a_495_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_207_n100# a_n705_n197# a_111_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_399_n100# a_n705_n197# a_303_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_495_n100# a_n705_n197# a_399_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_687_n100# a_n705_n197# a_591_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n561_n100# a_n705_n197# a_n657_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n465_n100# a_n705_n197# a_n561_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n657_n100# a_n705_n197# a_n749_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n369_n100# a_n705_n197# a_n465_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_15_n100# a_n705_n197# a_n81_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_111_n100# a_n705_n197# a_15_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n273_n100# a_n705_n197# a_n369_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n81_n100# a_n705_n197# a_n177_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n177_n100# a_n705_n197# a_n273_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_495_n100# a_687_n100# 0.11fF
C1 a_n749_n100# a_n369_n100# 0.05fF
C2 a_n657_n100# a_n705_n197# 0.08fF
C3 a_n81_n100# w_n887_n319# 0.02fF
C4 a_495_n100# w_n887_n319# 0.04fF
C5 a_n705_n197# a_n369_n100# 0.08fF
C6 a_15_n100# a_n177_n100# 0.11fF
C7 a_15_n100# w_n887_n319# 0.02fF
C8 a_495_n100# a_399_n100# 0.29fF
C9 a_n465_n100# a_n749_n100# 0.06fF
C10 a_n705_n197# a_n177_n100# 0.08fF
C11 a_111_n100# a_n273_n100# 0.05fF
C12 a_n465_n100# a_n705_n197# 0.08fF
C13 a_687_n100# a_303_n100# 0.05fF
C14 a_n749_n100# w_n887_n319# 0.10fF
C15 a_303_n100# w_n887_n319# 0.02fF
C16 a_n705_n197# w_n887_n319# 0.82fF
C17 a_n749_n100# a_n561_n100# 0.11fF
C18 a_687_n100# a_591_n100# 0.29fF
C19 a_15_n100# a_399_n100# 0.05fF
C20 a_591_n100# w_n887_n319# 0.05fF
C21 a_n705_n197# a_n561_n100# 0.08fF
C22 a_n81_n100# a_15_n100# 0.29fF
C23 a_399_n100# a_303_n100# 0.29fF
C24 a_n177_n100# a_111_n100# 0.06fF
C25 a_207_n100# a_n177_n100# 0.05fF
C26 a_n705_n197# a_399_n100# 0.08fF
C27 a_399_n100# a_591_n100# 0.11fF
C28 a_n81_n100# a_303_n100# 0.05fF
C29 a_495_n100# a_303_n100# 0.11fF
C30 a_n81_n100# a_n705_n197# 0.08fF
C31 a_n705_n197# a_495_n100# 0.08fF
C32 a_111_n100# w_n887_n319# 0.02fF
C33 a_207_n100# w_n887_n319# 0.02fF
C34 a_495_n100# a_591_n100# 0.29fF
C35 a_n657_n100# a_n273_n100# 0.05fF
C36 a_15_n100# a_303_n100# 0.06fF
C37 a_n369_n100# a_n273_n100# 0.29fF
C38 a_15_n100# a_n705_n197# 0.08fF
C39 a_399_n100# a_111_n100# 0.06fF
C40 a_n657_n100# a_n369_n100# 0.06fF
C41 a_207_n100# a_399_n100# 0.11fF
C42 a_n705_n197# a_303_n100# 0.08fF
C43 a_n81_n100# a_111_n100# 0.11fF
C44 a_495_n100# a_111_n100# 0.05fF
C45 a_n177_n100# a_n273_n100# 0.29fF
C46 a_207_n100# a_n81_n100# 0.06fF
C47 a_207_n100# a_495_n100# 0.06fF
C48 a_303_n100# a_591_n100# 0.06fF
C49 a_n465_n100# a_n273_n100# 0.11fF
C50 a_n705_n197# a_591_n100# 0.08fF
C51 a_n369_n100# a_n177_n100# 0.11fF
C52 a_n657_n100# a_n465_n100# 0.11fF
C53 a_n273_n100# w_n887_n319# 0.02fF
C54 a_15_n100# a_111_n100# 0.29fF
C55 a_207_n100# a_15_n100# 0.11fF
C56 a_n465_n100# a_n369_n100# 0.29fF
C57 a_n561_n100# a_n273_n100# 0.06fF
C58 a_n657_n100# w_n887_n319# 0.05fF
C59 a_n369_n100# w_n887_n319# 0.02fF
C60 a_n657_n100# a_n561_n100# 0.29fF
C61 a_303_n100# a_111_n100# 0.11fF
C62 a_207_n100# a_303_n100# 0.29fF
C63 a_n369_n100# a_n561_n100# 0.11fF
C64 a_n705_n197# a_111_n100# 0.08fF
C65 a_207_n100# a_n705_n197# 0.08fF
C66 a_n465_n100# a_n177_n100# 0.06fF
C67 a_207_n100# a_591_n100# 0.05fF
C68 a_n81_n100# a_n273_n100# 0.11fF
C69 a_n177_n100# w_n887_n319# 0.02fF
C70 a_n465_n100# w_n887_n319# 0.03fF
C71 a_n177_n100# a_n561_n100# 0.05fF
C72 a_687_n100# w_n887_n319# 0.10fF
C73 a_n81_n100# a_n369_n100# 0.06fF
C74 a_n465_n100# a_n561_n100# 0.29fF
C75 a_15_n100# a_n273_n100# 0.06fF
C76 a_n561_n100# w_n887_n319# 0.04fF
C77 a_207_n100# a_111_n100# 0.29fF
C78 a_15_n100# a_n369_n100# 0.05fF
C79 a_n81_n100# a_n177_n100# 0.29fF
C80 a_687_n100# a_399_n100# 0.06fF
C81 a_399_n100# w_n887_n319# 0.03fF
C82 a_n705_n197# a_n273_n100# 0.08fF
C83 a_n81_n100# a_n465_n100# 0.05fF
C84 a_n657_n100# a_n749_n100# 0.29fF
C85 a_687_n100# VSUBS 0.03fF
C86 a_591_n100# VSUBS 0.03fF
C87 a_495_n100# VSUBS 0.03fF
C88 a_399_n100# VSUBS 0.03fF
C89 a_303_n100# VSUBS 0.03fF
C90 a_207_n100# VSUBS 0.03fF
C91 a_111_n100# VSUBS 0.03fF
C92 a_15_n100# VSUBS 0.03fF
C93 a_n81_n100# VSUBS 0.03fF
C94 a_n177_n100# VSUBS 0.03fF
C95 a_n273_n100# VSUBS 0.03fF
C96 a_n369_n100# VSUBS 0.03fF
C97 a_n465_n100# VSUBS 0.03fF
C98 a_n561_n100# VSUBS 0.03fF
C99 a_n657_n100# VSUBS 0.03fF
C100 a_n749_n100# VSUBS 0.03fF
C101 a_n705_n197# VSUBS 1.60fF
C102 w_n887_n319# VSUBS 5.82fF
.ends

.subckt source_follower_buff_pmos m1_957_828# in avss1p8 avdd1p8 out iref
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_0 avss1p8 iref iref iref avss1p8 avss1p8 avss1p8
+ avss1p8 iref sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_1 avss1p8 m1_957_828# m1_957_828# iref avss1p8
+ avss1p8 avss1p8 avss1p8 m1_957_828# sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__pfet_01v8_lvt_D3F744_0 avss1p8 out avss1p8 out avss1p8 avss1p8 in out
+ avss1p8 avdd1p8 avss1p8 out out avss1p8 sky130_fd_pr__pfet_01v8_lvt_D3F744
Xsky130_fd_pr__pfet_01v8_VCU74W_0 avss1p8 m1_957_828# m1_957_828# avdd1p8 m1_957_828#
+ avdd1p8 m1_957_828# m1_957_828# avdd1p8 avdd1p8 avdd1p8 m1_957_828# m1_957_828#
+ m1_957_828# avdd1p8 avdd1p8 avdd1p8 m1_957_828# avdd1p8 sky130_fd_pr__pfet_01v8_VCU74W
Xsky130_fd_pr__pfet_01v8_VCU74W_1 avss1p8 out out avdd1p8 out avdd1p8 out out avdd1p8
+ avdd1p8 avdd1p8 out m1_957_828# out avdd1p8 avdd1p8 avdd1p8 out avdd1p8 sky130_fd_pr__pfet_01v8_VCU74W
C0 m1_957_828# avdd1p8 1.12fF
C1 in m1_957_828# 0.52fF
C2 m1_957_828# out 1.52fF
C3 m1_957_828# iref 0.88fF
C4 in avdd1p8 0.32fF
C5 avdd1p8 out 3.96fF
C6 iref avdd1p8 0.29fF
C7 in out 1.16fF
C8 avdd1p8 avss1p8 15.90fF
C9 out avss1p8 -1.64fF
C10 in avss1p8 1.94fF
C11 m1_957_828# avss1p8 -34.25fF
C12 iref avss1p8 4.22fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_CFLRKA a_n993_109# a_n1473_n309# a_63_n309# a_1215_n309#
+ a_1215_109# a_n129_n309# a_735_109# a_1599_109# a_n513_n309# a_255_109# a_n1377_n309#
+ a_n1949_109# a_n1761_n309# a_1119_n309# a_1503_n309# a_n1761_109# a_n417_109# a_n417_n309#
+ a_n1281_109# a_n801_n309# a_351_n309# a_63_109# a_1503_109# a_n1665_n309# a_1023_109#
+ a_1887_109# a_1407_n309# a_543_109# a_n705_n309# a_255_n309# a_1791_n309# a_n1569_109#
+ a_n705_109# a_n1569_n309# a_n1089_109# w_n2087_n519# a_n225_109# a_n609_n309# a_159_n309#
+ a_543_n309# a_1695_n309# a_1311_109# a_831_109# a_1695_109# a_n1857_n309# a_n993_n309#
+ a_n33_109# a_351_109# a_n1857_109# a_447_n309# a_831_n309# a_1599_n309# a_n1377_109#
+ a_n897_n309# a_n897_109# a_n513_109# a_1119_109# a_639_109# a_n33_n309# a_735_n309#
+ a_1887_n309# a_159_109# a_n1665_109# a_n1281_n309# a_1023_n309# a_n1185_109# a_n801_109#
+ a_639_n309# a_n321_109# a_1407_109# a_n321_n309# a_927_109# a_447_109# a_1791_109#
+ a_n1185_n309# a_1311_n309# a_n1905_n87# a_927_n309# a_n609_109# a_n225_n309# a_n1473_109#
+ a_n129_109# a_n1949_n309# a_n1089_n309#
X0 a_n1569_n309# a_n1905_n87# a_n1665_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n897_n309# a_n1905_n87# a_n993_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_927_n309# a_n1905_n87# a_831_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_1023_109# a_n1905_n87# a_927_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_255_n309# a_n1905_n87# a_159_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1215_n309# a_n1905_n87# a_1119_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_927_109# a_n1905_n87# a_831_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n1857_n309# a_n1905_n87# a_n1949_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n321_n309# a_n1905_n87# a_n417_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n1761_109# a_n1905_n87# a_n1857_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_543_n309# a_n1905_n87# a_447_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_1503_n309# a_n1905_n87# a_1407_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n1857_109# a_n1905_n87# a_n1949_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n1665_109# a_n1905_n87# a_n1761_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n1569_109# a_n1905_n87# a_n1665_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1215_109# a_n1905_n87# a_1119_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_1311_109# a_n1905_n87# a_1215_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_1503_109# a_n1905_n87# a_1407_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_1791_109# a_n1905_n87# a_1695_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n1185_n309# a_n1905_n87# a_n1281_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_1119_109# a_n1905_n87# a_1023_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1407_109# a_n1905_n87# a_1311_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1599_109# a_n1905_n87# a_1503_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_1695_109# a_n1905_n87# a_1599_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_1887_109# a_n1905_n87# a_1791_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_n1473_n309# a_n1905_n87# a_n1569_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_831_n309# a_n1905_n87# a_735_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_1791_n309# a_n1905_n87# a_1695_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n33_109# a_n1905_n87# a_n129_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_351_109# a_n1905_n87# a_255_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_159_n309# a_n1905_n87# a_63_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1119_n309# a_n1905_n87# a_1023_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_159_109# a_n1905_n87# a_63_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_255_109# a_n1905_n87# a_159_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_447_109# a_n1905_n87# a_351_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_543_109# a_n1905_n87# a_447_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_735_109# a_n1905_n87# a_639_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_831_109# a_n1905_n87# a_735_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n225_n309# a_n1905_n87# a_n321_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_639_109# a_n1905_n87# a_543_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_447_n309# a_n1905_n87# a_351_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_1407_n309# a_n1905_n87# a_1311_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_n1473_109# a_n1905_n87# a_n1569_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 a_n1281_109# a_n1905_n87# a_n1377_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 a_n1185_109# a_n1905_n87# a_n1281_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 a_n993_109# a_n1905_n87# a_n1089_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 a_n1089_n309# a_n1905_n87# a_n1185_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 a_n1377_109# a_n1905_n87# a_n1473_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_n1089_109# a_n1905_n87# a_n1185_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 a_n321_109# a_n1905_n87# a_n417_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n513_n309# a_n1905_n87# a_n609_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 a_63_n309# a_n1905_n87# a_n33_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_n801_109# a_n1905_n87# a_n897_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 a_n705_109# a_n1905_n87# a_n801_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_n513_109# a_n1905_n87# a_n609_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_n417_109# a_n1905_n87# a_n513_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 a_n225_109# a_n1905_n87# a_n321_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 a_n129_109# a_n1905_n87# a_n225_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_n1377_n309# a_n1905_n87# a_n1473_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 a_735_n309# a_n1905_n87# a_639_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X60 a_1695_n309# a_n1905_n87# a_1599_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 a_n897_109# a_n1905_n87# a_n993_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 a_n609_109# a_n1905_n87# a_n705_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 a_n801_n309# a_n1905_n87# a_n897_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 a_n129_n309# a_n1905_n87# a_n225_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 a_n1761_n309# a_n1905_n87# a_n1857_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 a_n417_n309# a_n1905_n87# a_n513_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 a_63_109# a_n1905_n87# a_n33_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 a_639_n309# a_n1905_n87# a_543_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 a_1599_n309# a_n1905_n87# a_1503_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 a_n705_n309# a_n1905_n87# a_n801_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X71 a_1887_n309# a_n1905_n87# a_1791_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 a_n1665_n309# a_n1905_n87# a_n1761_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 a_1023_n309# a_n1905_n87# a_927_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 a_n993_n309# a_n1905_n87# a_n1089_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 a_n33_n309# a_n1905_n87# a_n129_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 a_351_n309# a_n1905_n87# a_255_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 a_1311_n309# a_n1905_n87# a_1215_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 a_n1281_n309# a_n1905_n87# a_n1377_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X79 a_n609_n309# a_n1905_n87# a_n705_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_831_109# a_1119_109# 0.06fF
C1 a_n993_109# a_n1377_109# 0.05fF
C2 a_1887_n309# a_1695_n309# 0.11fF
C3 a_n897_109# a_n705_109# 0.11fF
C4 a_n417_n309# a_n129_n309# 0.06fF
C5 a_1503_109# a_1791_109# 0.06fF
C6 a_63_n309# a_n225_n309# 0.06fF
C7 a_1791_109# a_1599_109# 0.11fF
C8 a_831_109# a_447_109# 0.05fF
C9 a_n897_n309# a_n1089_n309# 0.11fF
C10 a_n417_109# a_n801_109# 0.05fF
C11 a_1023_n309# a_831_n309# 0.11fF
C12 a_n1857_n309# a_n1949_n309# 0.29fF
C13 a_n1569_n309# a_n1569_109# 0.01fF
C14 a_351_109# a_n33_109# 0.05fF
C15 a_639_109# a_1023_109# 0.05fF
C16 a_n1569_109# a_n1949_109# 0.05fF
C17 a_927_109# a_1215_109# 0.06fF
C18 a_63_n309# a_n321_n309# 0.05fF
C19 a_1023_n309# a_639_n309# 0.05fF
C20 a_159_n309# a_63_n309# 0.29fF
C21 a_n897_n309# a_n993_n309# 0.29fF
C22 a_n1281_n309# a_n1377_n309# 0.29fF
C23 a_n129_109# a_n225_109# 0.29fF
C24 a_n801_109# a_n897_109# 0.29fF
C25 a_1407_109# a_1023_109# 0.05fF
C26 a_n129_n309# a_255_n309# 0.05fF
C27 a_735_n309# a_1119_n309# 0.05fF
C28 a_63_109# a_n33_109# 0.29fF
C29 a_n1473_n309# a_n1089_n309# 0.05fF
C30 a_n897_n309# a_n1185_n309# 0.06fF
C31 a_351_n309# a_735_n309# 0.05fF
C32 a_n705_n309# a_n897_n309# 0.11fF
C33 a_63_109# a_n321_109# 0.05fF
C34 a_639_109# a_735_109# 0.29fF
C35 a_1503_109# a_1599_109# 0.29fF
C36 a_n993_109# a_n705_109# 0.06fF
C37 a_n129_109# a_255_109# 0.05fF
C38 a_831_109# a_1023_109# 0.11fF
C39 a_n705_n309# a_n321_n309# 0.05fF
C40 a_n1089_n309# a_n993_n309# 0.29fF
C41 a_159_109# a_n33_109# 0.11fF
C42 a_1119_n309# a_1503_n309# 0.05fF
C43 a_1215_n309# a_1503_n309# 0.06fF
C44 a_n1089_n309# a_n1185_n309# 0.29fF
C45 a_n801_n309# a_n417_n309# 0.05fF
C46 a_n1665_109# a_n1665_n309# 0.01fF
C47 a_447_n309# a_831_n309# 0.05fF
C48 a_n705_n309# a_n1089_n309# 0.05fF
C49 a_n225_n309# a_n513_n309# 0.06fF
C50 a_n417_109# a_n33_109# 0.05fF
C51 a_n1473_n309# a_n1185_n309# 0.06fF
C52 a_1119_109# a_1023_109# 0.29fF
C53 a_1503_109# a_1311_109# 0.11fF
C54 a_1599_109# a_1311_109# 0.06fF
C55 a_n417_109# a_n321_109# 0.29fF
C56 a_n1857_109# a_n1949_109# 0.29fF
C57 a_831_109# a_735_109# 0.29fF
C58 a_n897_n309# a_n513_n309# 0.05fF
C59 a_1791_n309# a_1599_n309# 0.11fF
C60 a_447_n309# a_639_n309# 0.11fF
C61 a_1887_109# a_1695_109# 0.11fF
C62 a_1311_n309# a_1599_n309# 0.06fF
C63 a_543_n309# a_831_n309# 0.06fF
C64 a_n993_109# a_n801_109# 0.11fF
C65 a_927_109# a_543_109# 0.05fF
C66 a_n993_n309# a_n1185_n309# 0.11fF
C67 a_n321_n309# a_n513_n309# 0.11fF
C68 a_n705_n309# a_n993_n309# 0.06fF
C69 a_1791_109# a_1791_n309# 0.01fF
C70 a_n1761_109# a_n1949_109# 0.11fF
C71 a_1119_109# a_735_109# 0.05fF
C72 a_1695_n309# a_1599_n309# 0.29fF
C73 a_n1761_n309# a_n1761_109# 0.01fF
C74 a_n801_109# a_n705_109# 0.29fF
C75 a_543_n309# a_639_n309# 0.29fF
C76 a_n417_109# a_n609_109# 0.11fF
C77 a_n129_109# a_n513_109# 0.05fF
C78 a_1023_n309# a_1407_n309# 0.05fF
C79 a_n1281_109# a_n1185_109# 0.29fF
C80 a_n897_n309# a_n1281_n309# 0.05fF
C81 a_543_109# a_351_109# 0.11fF
C82 a_n1089_109# a_n1089_n309# 0.01fF
C83 a_447_109# a_735_109# 0.06fF
C84 a_63_109# a_n225_109# 0.06fF
C85 a_n513_109# a_n513_n309# 0.01fF
C86 a_255_109# a_351_109# 0.29fF
C87 a_1215_109# a_1407_109# 0.11fF
C88 a_n1281_109# a_n1089_109# 0.11fF
C89 a_n1473_n309# a_n1473_109# 0.01fF
C90 a_n1185_109# a_n1185_n309# 0.01fF
C91 a_n897_109# a_n609_109# 0.06fF
C92 a_927_n309# a_1023_n309# 0.29fF
C93 a_n417_n309# a_n33_n309# 0.05fF
C94 a_1215_n309# a_1215_109# 0.01fF
C95 a_n1281_109# a_n1473_109# 0.11fF
C96 a_n1089_n309# a_n1281_n309# 0.11fF
C97 a_1791_n309# a_1407_n309# 0.05fF
C98 a_543_n309# a_543_109# 0.01fF
C99 a_63_109# a_255_109# 0.11fF
C100 a_n1473_n309# a_n1281_n309# 0.11fF
C101 a_1407_n309# a_1311_n309# 0.29fF
C102 a_159_109# a_n225_109# 0.05fF
C103 a_n1377_109# a_n1377_n309# 0.01fF
C104 a_639_109# a_639_n309# 0.01fF
C105 a_831_109# a_1215_109# 0.05fF
C106 a_n1665_109# a_n1949_109# 0.06fF
C107 a_n1281_109# a_n1281_n309# 0.01fF
C108 a_n801_n309# a_n609_n309# 0.11fF
C109 a_n705_n309# a_n513_n309# 0.11fF
C110 a_831_n309# a_1119_n309# 0.06fF
C111 a_1215_n309# a_831_n309# 0.05fF
C112 a_159_109# a_543_109# 0.05fF
C113 a_n417_109# a_n225_109# 0.11fF
C114 a_1695_n309# a_1407_n309# 0.06fF
C115 a_255_n309# a_639_n309# 0.05fF
C116 a_1791_109# a_1695_109# 0.29fF
C117 a_n1857_109# a_n1857_n309# 0.01fF
C118 a_159_n309# a_447_n309# 0.06fF
C119 a_n993_n309# a_n1281_n309# 0.06fF
C120 a_735_109# a_735_n309# 0.01fF
C121 a_n417_n309# a_n225_n309# 0.11fF
C122 a_1215_109# a_1119_109# 0.29fF
C123 a_159_109# a_255_109# 0.29fF
C124 a_927_n309# a_927_109# 0.01fF
C125 a_735_109# a_1023_109# 0.06fF
C126 a_831_109# a_831_n309# 0.01fF
C127 a_n609_n309# a_n609_109# 0.01fF
C128 a_n33_n309# a_255_n309# 0.06fF
C129 a_n1281_n309# a_n1185_n309# 0.29fF
C130 a_927_n309# a_1311_n309# 0.05fF
C131 a_n1281_109# a_n1569_109# 0.06fF
C132 a_351_n309# a_639_n309# 0.06fF
C133 a_447_n309# a_63_n309# 0.05fF
C134 a_n1185_109# a_n1089_109# 0.29fF
C135 a_n321_109# a_n705_109# 0.05fF
C136 a_927_109# a_1311_109# 0.05fF
C137 a_159_n309# a_543_n309# 0.05fF
C138 a_639_109# a_543_109# 0.29fF
C139 a_n1185_109# a_n1473_109# 0.06fF
C140 a_1311_109# a_1311_n309# 0.01fF
C141 a_63_n309# a_63_109# 0.01fF
C142 a_n417_n309# a_n321_n309# 0.29fF
C143 a_n33_n309# a_351_n309# 0.05fF
C144 a_639_109# a_255_109# 0.05fF
C145 a_n993_109# a_n609_109# 0.05fF
C146 a_159_n309# a_159_109# 0.01fF
C147 a_1215_n309# a_1599_n309# 0.05fF
C148 a_n1569_n309# a_n1665_n309# 0.29fF
C149 a_255_109# a_255_n309# 0.01fF
C150 a_1791_109# a_1407_109# 0.05fF
C151 a_n705_109# a_n609_109# 0.29fF
C152 a_n1089_109# a_n1473_109# 0.05fF
C153 a_n1761_n309# a_n1665_n309# 0.29fF
C154 a_1503_109# a_1695_109# 0.11fF
C155 a_1599_109# a_1695_109# 0.29fF
C156 a_1887_n309# a_1503_n309# 0.05fF
C157 a_927_n309# a_543_n309# 0.05fF
C158 a_n897_n309# a_n897_109# 0.01fF
C159 a_831_109# a_543_109# 0.06fF
C160 a_n801_n309# a_n801_109# 0.01fF
C161 a_n1185_109# a_n1569_109# 0.05fF
C162 a_1023_n309# a_1311_n309# 0.06fF
C163 a_n417_109# a_n513_109# 0.29fF
C164 a_159_n309# a_255_n309# 0.29fF
C165 a_1215_109# a_1023_109# 0.11fF
C166 a_1311_109# a_1695_109# 0.05fF
C167 a_n801_109# a_n609_109# 0.11fF
C168 a_n1665_n309# a_n1377_n309# 0.06fF
C169 a_1407_n309# a_1407_109# 0.01fF
C170 a_n705_n309# a_n417_n309# 0.06fF
C171 a_n129_109# a_63_109# 0.11fF
C172 a_n225_n309# a_n609_n309# 0.05fF
C173 a_63_n309# a_255_n309# 0.11fF
C174 a_1407_n309# a_1119_n309# 0.06fF
C175 a_159_n309# a_351_n309# 0.11fF
C176 a_735_n309# a_831_n309# 0.29fF
C177 a_447_109# a_543_109# 0.29fF
C178 a_n1473_109# a_n1569_109# 0.29fF
C179 a_1215_n309# a_1407_n309# 0.11fF
C180 a_1503_109# a_1407_109# 0.29fF
C181 a_n897_n309# a_n609_n309# 0.06fF
C182 a_1599_109# a_1407_109# 0.11fF
C183 a_n513_109# a_n897_109# 0.05fF
C184 a_n1281_109# a_n897_109# 0.05fF
C185 a_447_109# a_255_109# 0.11fF
C186 a_63_n309# a_351_n309# 0.06fF
C187 a_735_n309# a_639_n309# 0.29fF
C188 a_n1377_109# a_n1281_109# 0.29fF
C189 a_n321_n309# a_n609_n309# 0.06fF
C190 a_1791_n309# a_1695_n309# 0.29fF
C191 a_n129_109# a_159_109# 0.06fF
C192 a_1695_n309# a_1311_n309# 0.05fF
C193 a_927_n309# a_1119_n309# 0.11fF
C194 a_n1761_n309# a_n1569_n309# 0.11fF
C195 a_n417_109# a_n129_109# 0.06fF
C196 a_1215_n309# a_927_n309# 0.06fF
C197 a_1311_109# a_1407_109# 0.29fF
C198 a_n417_n309# a_n513_n309# 0.29fF
C199 a_n321_109# a_n33_109# 0.06fF
C200 a_n1857_n309# a_n1665_n309# 0.11fF
C201 a_1887_n309# a_1887_109# 0.01fF
C202 a_n33_n309# a_n129_n309# 0.29fF
C203 a_1503_109# a_1119_109# 0.05fF
C204 a_n1281_109# a_n1665_109# 0.05fF
C205 a_n1185_109# a_n897_109# 0.06fF
C206 a_n993_n309# a_n609_n309# 0.05fF
C207 a_n1569_n309# a_n1377_n309# 0.11fF
C208 a_63_109# a_351_109# 0.06fF
C209 a_n1857_109# a_n1473_109# 0.05fF
C210 a_n1377_109# a_n1185_109# 0.11fF
C211 a_n321_109# a_n609_109# 0.06fF
C212 a_n993_109# a_n1281_109# 0.06fF
C213 a_1503_n309# a_1599_n309# 0.29fF
C214 a_n129_n309# a_n225_n309# 0.29fF
C215 a_n1761_n309# a_n1377_n309# 0.05fF
C216 a_n705_n309# a_n609_n309# 0.29fF
C217 a_1311_109# a_1119_109# 0.11fF
C218 a_447_n309# a_543_n309# 0.29fF
C219 a_n1089_109# a_n897_109# 0.11fF
C220 a_n513_109# a_n705_109# 0.11fF
C221 a_1023_n309# a_1119_n309# 0.29fF
C222 a_1695_n309# a_1695_109# 0.01fF
C223 a_n993_109# a_n993_n309# 0.01fF
C224 a_n1761_109# a_n1473_109# 0.06fF
C225 a_543_109# a_735_109# 0.11fF
C226 a_1215_n309# a_1023_n309# 0.11fF
C227 a_n1377_109# a_n1089_109# 0.06fF
C228 a_159_109# a_351_109# 0.11fF
C229 a_639_109# a_927_109# 0.06fF
C230 a_n1377_109# a_n1473_109# 0.29fF
C231 a_n321_n309# a_n129_n309# 0.11fF
C232 a_1887_n309# a_1599_n309# 0.06fF
C233 a_159_n309# a_n129_n309# 0.06fF
C234 a_n33_n309# a_n33_109# 0.01fF
C235 a_n1857_109# a_n1569_109# 0.06fF
C236 a_n1473_n309# a_n1665_n309# 0.11fF
C237 a_n1569_n309# a_n1857_n309# 0.06fF
C238 a_n705_n309# a_n705_109# 0.01fF
C239 a_159_109# a_63_109# 0.29fF
C240 a_n225_109# a_n33_109# 0.11fF
C241 a_639_109# a_351_109# 0.06fF
C242 a_n513_n309# a_n609_n309# 0.29fF
C243 a_63_n309# a_n129_n309# 0.11fF
C244 a_n801_109# a_n513_109# 0.06fF
C245 a_n1761_n309# a_n1857_n309# 0.29fF
C246 a_n993_109# a_n1185_109# 0.11fF
C247 a_n225_109# a_n321_109# 0.29fF
C248 a_1311_n309# a_1119_n309# 0.11fF
C249 a_n1761_109# a_n1569_109# 0.11fF
C250 a_1215_n309# a_1311_n309# 0.29fF
C251 a_927_n309# a_735_n309# 0.11fF
C252 a_1407_n309# a_1503_n309# 0.29fF
C253 a_831_109# a_927_109# 0.29fF
C254 a_447_n309# a_255_n309# 0.11fF
C255 a_n1665_109# a_n1473_109# 0.11fF
C256 a_n1377_109# a_n1569_109# 0.11fF
C257 a_255_109# a_n33_109# 0.06fF
C258 a_831_n309# a_639_n309# 0.11fF
C259 a_n993_109# a_n1089_109# 0.29fF
C260 a_1503_109# a_1503_n309# 0.01fF
C261 a_n1665_n309# a_n1949_n309# 0.06fF
C262 a_351_n309# a_351_109# 0.01fF
C263 a_n417_109# a_n417_n309# 0.01fF
C264 a_1311_109# a_1023_109# 0.06fF
C265 a_n225_109# a_n609_109# 0.05fF
C266 a_447_n309# a_351_n309# 0.29fF
C267 a_927_109# a_1119_109# 0.11fF
C268 a_n1089_109# a_n705_109# 0.05fF
C269 a_543_n309# a_255_n309# 0.06fF
C270 a_n897_n309# a_n801_n309# 0.29fF
C271 a_1791_109# a_1887_109# 0.29fF
C272 a_n321_n309# a_n321_109# 0.01fF
C273 a_1407_109# a_1695_109# 0.06fF
C274 a_n801_109# a_n1185_109# 0.05fF
C275 a_543_n309# a_351_n309# 0.11fF
C276 a_n1665_109# a_n1569_109# 0.29fF
C277 a_n129_109# a_n129_n309# 0.01fF
C278 a_n1569_n309# a_n1473_n309# 0.29fF
C279 a_1023_n309# a_735_n309# 0.06fF
C280 a_n1857_109# a_n1761_109# 0.29fF
C281 a_1023_n309# a_1023_109# 0.01fF
C282 a_447_109# a_351_109# 0.29fF
C283 a_n801_n309# a_n1089_n309# 0.06fF
C284 a_n801_109# a_n1089_109# 0.06fF
C285 a_n1761_n309# a_n1473_n309# 0.06fF
C286 a_n129_n309# a_n513_n309# 0.05fF
C287 a_447_n309# a_447_109# 0.01fF
C288 a_n513_109# a_n321_109# 0.11fF
C289 a_447_109# a_63_109# 0.05fF
C290 a_n1665_n309# a_n1281_n309# 0.05fF
C291 a_n1569_n309# a_n1185_n309# 0.05fF
C292 a_1503_109# a_1215_109# 0.06fF
C293 a_n417_n309# a_n609_n309# 0.11fF
C294 a_1599_109# a_1215_109# 0.05fF
C295 a_n1569_n309# a_n1949_n309# 0.05fF
C296 a_n801_n309# a_n993_n309# 0.11fF
C297 a_n33_n309# a_n225_n309# 0.11fF
C298 a_n1089_n309# a_n1377_n309# 0.06fF
C299 a_n1377_109# a_n1761_109# 0.05fF
C300 a_1503_109# a_1887_109# 0.05fF
C301 a_1599_109# a_1887_109# 0.06fF
C302 a_927_109# a_1023_109# 0.29fF
C303 a_n513_109# a_n609_109# 0.29fF
C304 a_n1949_109# a_n1949_n309# 0.01fF
C305 a_831_109# a_639_109# 0.11fF
C306 a_n1473_n309# a_n1377_n309# 0.29fF
C307 a_n225_n309# a_n225_109# 0.01fF
C308 a_351_n309# a_255_n309# 0.29fF
C309 a_n1761_n309# a_n1949_n309# 0.11fF
C310 a_n801_n309# a_n1185_n309# 0.05fF
C311 a_n705_n309# a_n801_n309# 0.29fF
C312 a_1215_n309# a_1119_n309# 0.29fF
C313 a_159_109# a_447_109# 0.06fF
C314 a_543_109# a_255_109# 0.06fF
C315 a_n1857_109# a_n1665_109# 0.11fF
C316 a_n33_n309# a_n321_n309# 0.06fF
C317 a_1215_109# a_1311_109# 0.29fF
C318 a_n129_109# a_n33_109# 0.29fF
C319 a_n993_n309# a_n1377_n309# 0.05fF
C320 a_447_n309# a_735_n309# 0.06fF
C321 a_1791_n309# a_1503_n309# 0.06fF
C322 a_159_n309# a_n33_n309# 0.11fF
C323 a_n129_109# a_n321_109# 0.11fF
C324 a_927_109# a_735_109# 0.11fF
C325 a_927_n309# a_831_n309# 0.29fF
C326 a_1311_n309# a_1503_n309# 0.11fF
C327 a_n1377_n309# a_n1185_n309# 0.11fF
C328 a_n1761_109# a_n1665_109# 0.29fF
C329 a_1119_109# a_1407_109# 0.06fF
C330 a_639_109# a_447_109# 0.11fF
C331 a_n33_n309# a_63_n309# 0.29fF
C332 a_n417_109# a_n705_109# 0.06fF
C333 a_1407_n309# a_1599_n309# 0.11fF
C334 a_1695_n309# a_1503_n309# 0.11fF
C335 a_543_n309# a_735_n309# 0.11fF
C336 a_1119_109# a_1119_n309# 0.01fF
C337 a_927_n309# a_639_n309# 0.06fF
C338 a_n1377_109# a_n1665_109# 0.06fF
C339 a_n1473_n309# a_n1857_n309# 0.05fF
C340 a_735_109# a_351_109# 0.05fF
C341 a_1887_n309# a_1791_n309# 0.29fF
C342 a_n801_n309# a_n513_n309# 0.06fF
C343 a_n321_n309# a_n225_n309# 0.29fF
C344 a_n225_109# a_n513_109# 0.06fF
C345 a_n993_109# a_n897_109# 0.29fF
C346 a_159_n309# a_n225_n309# 0.05fF
C347 a_1599_109# a_1599_n309# 0.01fF
C348 a_n1569_n309# a_n1281_n309# 0.06fF
C349 a_1887_n309# w_n2087_n519# 0.12fF
C350 a_1791_n309# w_n2087_n519# 0.08fF
C351 a_1695_n309# w_n2087_n519# 0.06fF
C352 a_1599_n309# w_n2087_n519# 0.06fF
C353 a_1503_n309# w_n2087_n519# 0.04fF
C354 a_1407_n309# w_n2087_n519# 0.04fF
C355 a_1311_n309# w_n2087_n519# 0.04fF
C356 a_1215_n309# w_n2087_n519# 0.04fF
C357 a_1119_n309# w_n2087_n519# 0.04fF
C358 a_1023_n309# w_n2087_n519# 0.04fF
C359 a_927_n309# w_n2087_n519# 0.04fF
C360 a_831_n309# w_n2087_n519# 0.04fF
C361 a_735_n309# w_n2087_n519# 0.04fF
C362 a_639_n309# w_n2087_n519# 0.04fF
C363 a_543_n309# w_n2087_n519# 0.04fF
C364 a_447_n309# w_n2087_n519# 0.04fF
C365 a_351_n309# w_n2087_n519# 0.04fF
C366 a_255_n309# w_n2087_n519# 0.04fF
C367 a_159_n309# w_n2087_n519# 0.04fF
C368 a_63_n309# w_n2087_n519# 0.04fF
C369 a_n33_n309# w_n2087_n519# 0.04fF
C370 a_n129_n309# w_n2087_n519# 0.04fF
C371 a_n225_n309# w_n2087_n519# 0.04fF
C372 a_n321_n309# w_n2087_n519# 0.04fF
C373 a_n417_n309# w_n2087_n519# 0.04fF
C374 a_n513_n309# w_n2087_n519# 0.04fF
C375 a_n609_n309# w_n2087_n519# 0.04fF
C376 a_n705_n309# w_n2087_n519# 0.04fF
C377 a_n801_n309# w_n2087_n519# 0.04fF
C378 a_n897_n309# w_n2087_n519# 0.04fF
C379 a_n993_n309# w_n2087_n519# 0.04fF
C380 a_n1089_n309# w_n2087_n519# 0.04fF
C381 a_n1185_n309# w_n2087_n519# 0.04fF
C382 a_n1281_n309# w_n2087_n519# 0.04fF
C383 a_n1377_n309# w_n2087_n519# 0.04fF
C384 a_n1473_n309# w_n2087_n519# 0.04fF
C385 a_n1569_n309# w_n2087_n519# 0.04fF
C386 a_n1665_n309# w_n2087_n519# 0.04fF
C387 a_n1761_n309# w_n2087_n519# 0.04fF
C388 a_n1857_n309# w_n2087_n519# 0.04fF
C389 a_n1949_n309# w_n2087_n519# 0.04fF
C390 a_1887_109# w_n2087_n519# 0.12fF
C391 a_1791_109# w_n2087_n519# 0.08fF
C392 a_1695_109# w_n2087_n519# 0.06fF
C393 a_1599_109# w_n2087_n519# 0.06fF
C394 a_1503_109# w_n2087_n519# 0.04fF
C395 a_1407_109# w_n2087_n519# 0.04fF
C396 a_1311_109# w_n2087_n519# 0.04fF
C397 a_1215_109# w_n2087_n519# 0.04fF
C398 a_1119_109# w_n2087_n519# 0.04fF
C399 a_1023_109# w_n2087_n519# 0.04fF
C400 a_927_109# w_n2087_n519# 0.04fF
C401 a_831_109# w_n2087_n519# 0.04fF
C402 a_735_109# w_n2087_n519# 0.04fF
C403 a_639_109# w_n2087_n519# 0.04fF
C404 a_543_109# w_n2087_n519# 0.04fF
C405 a_447_109# w_n2087_n519# 0.04fF
C406 a_351_109# w_n2087_n519# 0.04fF
C407 a_255_109# w_n2087_n519# 0.04fF
C408 a_159_109# w_n2087_n519# 0.04fF
C409 a_63_109# w_n2087_n519# 0.04fF
C410 a_n33_109# w_n2087_n519# 0.04fF
C411 a_n129_109# w_n2087_n519# 0.04fF
C412 a_n225_109# w_n2087_n519# 0.04fF
C413 a_n321_109# w_n2087_n519# 0.04fF
C414 a_n417_109# w_n2087_n519# 0.04fF
C415 a_n513_109# w_n2087_n519# 0.04fF
C416 a_n609_109# w_n2087_n519# 0.04fF
C417 a_n705_109# w_n2087_n519# 0.04fF
C418 a_n801_109# w_n2087_n519# 0.04fF
C419 a_n897_109# w_n2087_n519# 0.04fF
C420 a_n993_109# w_n2087_n519# 0.04fF
C421 a_n1089_109# w_n2087_n519# 0.04fF
C422 a_n1185_109# w_n2087_n519# 0.04fF
C423 a_n1281_109# w_n2087_n519# 0.04fF
C424 a_n1377_109# w_n2087_n519# 0.04fF
C425 a_n1473_109# w_n2087_n519# 0.04fF
C426 a_n1569_109# w_n2087_n519# 0.04fF
C427 a_n1665_109# w_n2087_n519# 0.04fF
C428 a_n1761_109# w_n2087_n519# 0.04fF
C429 a_n1857_109# w_n2087_n519# 0.04fF
C430 a_n1949_109# w_n2087_n519# 0.04fF
C431 a_n1905_n87# w_n2087_n519# 6.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_CAF2P9 a_63_n309# a_n1473_n309# a_159_527# a_1215_n309#
+ a_n993_109# a_1215_109# a_n129_n309# a_n513_n309# a_1599_109# a_735_109# a_n1665_527#
+ a_n1281_n727# a_n801_527# a_1023_n727# a_639_n727# a_255_109# a_n1185_527# a_n1377_n309#
+ a_n1949_109# a_1119_n309# a_n1761_n309# a_n321_527# a_1503_n309# a_1407_527# a_n321_n727#
+ a_927_527# a_n1761_109# a_n417_109# a_n417_n309# a_351_n309# a_n801_n309# a_n1905_n505#
+ a_n1281_109# a_n1185_n727# a_447_527# a_1791_527# a_63_109# a_1311_n727# a_927_n727#
+ a_1503_109# a_n1665_n309# a_1407_n309# a_1887_109# a_n225_n727# a_1023_109# a_n609_527#
+ a_543_109# a_255_n309# a_n1473_527# a_n1949_n727# a_1791_n309# a_n705_n309# a_n129_527#
+ a_n1089_n727# a_n1473_n727# a_1215_n727# a_63_n727# a_n993_527# a_n1569_109# a_n1569_n309#
+ a_n705_109# a_1215_527# a_n129_n727# a_n1089_109# a_1599_527# a_n513_n727# a_735_527#
+ a_n225_109# a_1695_n309# a_159_n309# a_n609_n309# a_543_n309# a_255_527# a_n1377_n727#
+ a_n1949_527# a_1119_n727# a_n1761_n727# a_1503_n727# a_1311_109# a_n993_n309# a_1695_109#
+ a_n1857_n309# a_831_109# a_n1761_527# a_n33_109# a_n417_n727# a_n417_527# a_351_109#
+ a_351_n727# a_n801_n727# a_n1281_527# a_n1857_109# a_1599_n309# a_447_n309# a_63_527#
+ a_831_n309# a_1503_527# a_n1377_109# a_n1665_n727# a_1887_527# a_1407_n727# a_n897_n309#
+ a_1023_527# a_n513_109# a_n897_109# a_543_527# a_1791_n727# a_255_n727# a_n705_n727#
+ a_1119_109# a_1887_n309# a_639_109# a_735_n309# a_n33_n309# a_n1569_527# a_n1569_n727#
+ a_n705_527# a_159_109# a_n1089_527# a_n225_527# w_n2087_n937# a_1695_n727# a_159_n727#
+ a_n609_n727# a_543_n727# a_n1665_109# a_n1281_n309# a_1023_n309# a_1311_527# a_n801_109#
+ a_639_n309# a_1695_527# a_n1185_109# a_n993_n727# a_831_527# a_n1857_n727# a_n321_109#
+ a_1407_109# a_n33_527# a_n321_n309# a_351_527# a_927_109# a_1599_n727# a_n1857_527#
+ a_447_n727# a_831_n727# a_447_109# a_n1185_n309# a_n1377_527# a_1791_109# a_1311_n309#
+ a_n897_n727# a_927_n309# a_n513_527# a_n897_527# a_n225_n309# a_n609_109# a_1119_527#
+ a_1887_n727# a_n1949_n309# a_639_527# a_n1473_109# a_n129_109# a_735_n727# a_n33_n727#
+ a_n1089_n309#
X0 a_927_n309# a_n1905_n505# a_831_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n897_n309# a_n1905_n505# a_n993_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n1569_n309# a_n1905_n505# a_n1665_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n129_n727# a_n1905_n505# a_n225_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n1761_n727# a_n1905_n505# a_n1857_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1215_n309# a_n1905_n505# a_1119_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_255_n309# a_n1905_n505# a_159_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_1023_109# a_n1905_n505# a_927_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n1857_n309# a_n1905_n505# a_n1949_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_927_109# a_n1905_n505# a_831_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n417_n727# a_n1905_n505# a_n513_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n321_n309# a_n1905_n505# a_n417_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_1599_n727# a_n1905_n505# a_1503_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_63_527# a_n1905_n505# a_n33_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n1761_109# a_n1905_n505# a_n1857_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1503_n309# a_n1905_n505# a_1407_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_639_n727# a_n1905_n505# a_543_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_543_n309# a_n1905_n505# a_447_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n1665_109# a_n1905_n505# a_n1761_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n1185_n309# a_n1905_n505# a_n1281_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_n1569_109# a_n1905_n505# a_n1665_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1311_109# a_n1905_n505# a_1215_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_n1857_109# a_n1905_n505# a_n1949_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_1791_109# a_n1905_n505# a_1695_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_1503_109# a_n1905_n505# a_1407_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_1215_109# a_n1905_n505# a_1119_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_n705_n727# a_n1905_n505# a_n801_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_1119_109# a_n1905_n505# a_1023_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1695_109# a_n1905_n505# a_1599_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1407_109# a_n1905_n505# a_1311_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_1599_109# a_n1905_n505# a_1503_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1887_109# a_n1905_n505# a_1791_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1887_n727# a_n1905_n505# a_1791_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_1791_n309# a_n1905_n505# a_1695_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_831_n309# a_n1905_n505# a_735_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_n1473_n309# a_n1905_n505# a_n1569_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_n33_109# a_n1905_n505# a_n129_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_1023_n727# a_n1905_n505# a_927_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n1665_n727# a_n1905_n505# a_n1761_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_1119_n309# a_n1905_n505# a_1023_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_159_n309# a_n1905_n505# a_63_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_351_109# a_n1905_n505# a_255_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_1311_n727# a_n1905_n505# a_1215_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 a_255_109# a_n1905_n505# a_159_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 a_351_n727# a_n1905_n505# a_255_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 a_831_109# a_n1905_n505# a_735_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 a_543_109# a_n1905_n505# a_447_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 a_n33_n727# a_n1905_n505# a_n129_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_n993_n727# a_n1905_n505# a_n1089_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 a_159_109# a_n1905_n505# a_63_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n225_n309# a_n1905_n505# a_n321_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 a_735_109# a_n1905_n505# a_639_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_447_109# a_n1905_n505# a_351_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 a_639_109# a_n1905_n505# a_543_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_1407_n309# a_n1905_n505# a_1311_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_447_n309# a_n1905_n505# a_351_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 a_n1089_n309# a_n1905_n505# a_n1185_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 a_n1281_109# a_n1905_n505# a_n1377_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_n993_109# a_n1905_n505# a_n1089_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 a_n1473_109# a_n1905_n505# a_n1569_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X60 a_n1185_109# a_n1905_n505# a_n1281_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 a_n609_n727# a_n1905_n505# a_n705_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 a_n1377_109# a_n1905_n505# a_n1473_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 a_n1089_109# a_n1905_n505# a_n1185_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 a_n1281_n727# a_n1905_n505# a_n1377_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 a_n513_n309# a_n1905_n505# a_n609_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 a_n321_109# a_n1905_n505# a_n417_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 a_63_n309# a_n1905_n505# a_n33_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 a_n225_109# a_n1905_n505# a_n321_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 a_n801_109# a_n1905_n505# a_n897_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 a_n513_109# a_n1905_n505# a_n609_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X71 a_1695_n309# a_n1905_n505# a_1599_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 a_n705_109# a_n1905_n505# a_n801_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 a_n417_109# a_n1905_n505# a_n513_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 a_n129_109# a_n1905_n505# a_n225_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 a_735_n309# a_n1905_n505# a_639_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 a_n1377_n309# a_n1905_n505# a_n1473_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 a_n897_109# a_n1905_n505# a_n993_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 a_n609_109# a_n1905_n505# a_n705_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X79 a_927_n727# a_n1905_n505# a_831_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X80 a_n1569_n727# a_n1905_n505# a_n1665_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X81 a_n897_n727# a_n1905_n505# a_n993_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X82 a_n801_n309# a_n1905_n505# a_n897_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 a_1215_n727# a_n1905_n505# a_1119_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X84 a_255_n727# a_n1905_n505# a_159_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X85 a_1023_527# a_n1905_n505# a_927_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X86 a_n129_n309# a_n1905_n505# a_n225_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X87 a_927_527# a_n1905_n505# a_831_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X88 a_n1857_n727# a_n1905_n505# a_n1949_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X89 a_n1761_n309# a_n1905_n505# a_n1857_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X90 a_n321_n727# a_n1905_n505# a_n417_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X91 a_n1761_527# a_n1905_n505# a_n1857_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 a_1503_n727# a_n1905_n505# a_1407_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X93 a_n1665_527# a_n1905_n505# a_n1761_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X94 a_543_n727# a_n1905_n505# a_447_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X95 a_n1185_n727# a_n1905_n505# a_n1281_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X96 a_n417_n309# a_n1905_n505# a_n513_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X97 a_n1857_527# a_n1905_n505# a_n1949_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X98 a_n1569_527# a_n1905_n505# a_n1665_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 a_1311_527# a_n1905_n505# a_1215_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X100 a_1215_527# a_n1905_n505# a_1119_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 a_1503_527# a_n1905_n505# a_1407_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X102 a_1791_527# a_n1905_n505# a_1695_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X103 a_1119_527# a_n1905_n505# a_1023_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X104 a_1407_527# a_n1905_n505# a_1311_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X105 a_1695_527# a_n1905_n505# a_1599_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X106 a_1599_n309# a_n1905_n505# a_1503_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X107 a_63_109# a_n1905_n505# a_n33_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X108 a_639_n309# a_n1905_n505# a_543_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X109 a_1599_527# a_n1905_n505# a_1503_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X110 a_1887_527# a_n1905_n505# a_1791_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X111 a_1791_n727# a_n1905_n505# a_1695_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X112 a_831_n727# a_n1905_n505# a_735_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X113 a_n1473_n727# a_n1905_n505# a_n1569_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 a_n705_n309# a_n1905_n505# a_n801_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 a_n33_527# a_n1905_n505# a_n129_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 a_1887_n309# a_n1905_n505# a_1791_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X117 a_1119_n727# a_n1905_n505# a_1023_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 a_159_n727# a_n1905_n505# a_63_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X119 a_351_527# a_n1905_n505# a_255_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X120 a_1023_n309# a_n1905_n505# a_927_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X121 a_n1665_n309# a_n1905_n505# a_n1761_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X122 a_255_527# a_n1905_n505# a_159_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X123 a_543_527# a_n1905_n505# a_447_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X124 a_831_527# a_n1905_n505# a_735_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X125 a_159_527# a_n1905_n505# a_63_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X126 a_447_527# a_n1905_n505# a_351_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X127 a_n225_n727# a_n1905_n505# a_n321_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X128 a_735_527# a_n1905_n505# a_639_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X129 a_639_527# a_n1905_n505# a_543_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X130 a_1407_n727# a_n1905_n505# a_1311_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X131 a_447_n727# a_n1905_n505# a_351_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X132 a_1311_n309# a_n1905_n505# a_1215_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X133 a_n1089_n727# a_n1905_n505# a_n1185_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X134 a_351_n309# a_n1905_n505# a_255_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 a_n33_n309# a_n1905_n505# a_n129_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X136 a_n1281_527# a_n1905_n505# a_n1377_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X137 a_n993_527# a_n1905_n505# a_n1089_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X138 a_n993_n309# a_n1905_n505# a_n1089_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X139 a_n1473_527# a_n1905_n505# a_n1569_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 a_n1185_527# a_n1905_n505# a_n1281_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X141 a_n1377_527# a_n1905_n505# a_n1473_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X142 a_n1089_527# a_n1905_n505# a_n1185_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X143 a_n513_n727# a_n1905_n505# a_n609_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X144 a_n321_527# a_n1905_n505# a_n417_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X145 a_63_n727# a_n1905_n505# a_n33_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X146 a_n801_527# a_n1905_n505# a_n897_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X147 a_n513_527# a_n1905_n505# a_n609_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X148 a_n225_527# a_n1905_n505# a_n321_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X149 a_1695_n727# a_n1905_n505# a_1599_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X150 a_735_n727# a_n1905_n505# a_639_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X151 a_n705_527# a_n1905_n505# a_n801_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X152 a_n417_527# a_n1905_n505# a_n513_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X153 a_n129_527# a_n1905_n505# a_n225_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X154 a_n1377_n727# a_n1905_n505# a_n1473_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 a_n609_n309# a_n1905_n505# a_n705_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 a_n1281_n309# a_n1905_n505# a_n1377_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X157 a_n897_527# a_n1905_n505# a_n993_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X158 a_n609_527# a_n1905_n505# a_n705_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X159 a_n801_n727# a_n1905_n505# a_n897_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_735_n727# a_735_n309# 0.01fF
C1 a_n897_527# a_n1185_527# 0.06fF
C2 a_n1377_109# a_n1377_n309# 0.01fF
C3 a_n1665_n727# a_n1761_n727# 0.29fF
C4 a_255_109# a_159_109# 0.29fF
C5 a_1215_109# a_927_109# 0.06fF
C6 a_n225_n727# a_n225_n309# 0.01fF
C7 a_927_n727# a_1311_n727# 0.05fF
C8 a_n1949_527# a_n1569_527# 0.05fF
C9 a_831_527# a_1023_527# 0.11fF
C10 a_831_109# a_927_109# 0.29fF
C11 a_n705_109# a_n801_109# 0.29fF
C12 a_n33_527# a_n33_109# 0.01fF
C13 a_543_109# a_447_109# 0.29fF
C14 a_159_n309# a_447_n309# 0.06fF
C15 a_1023_n727# a_1215_n727# 0.11fF
C16 a_927_109# a_1023_109# 0.29fF
C17 a_1503_n309# a_1407_n309# 0.29fF
C18 a_n321_109# a_n225_109# 0.29fF
C19 a_543_n309# a_927_n309# 0.05fF
C20 a_n417_527# a_n129_527# 0.06fF
C21 a_n321_527# a_n33_527# 0.06fF
C22 a_831_n727# a_543_n727# 0.06fF
C23 a_639_n309# a_543_n309# 0.29fF
C24 a_n1185_n727# a_n897_n727# 0.06fF
C25 a_n321_n727# a_n705_n727# 0.05fF
C26 a_1311_n727# a_1215_n727# 0.29fF
C27 a_n1089_n727# a_n897_n727# 0.11fF
C28 a_n1281_527# a_n1569_527# 0.06fF
C29 a_1215_n309# a_1023_n309# 0.11fF
C30 a_n417_n309# a_n417_n727# 0.01fF
C31 a_n1377_527# a_n993_527# 0.05fF
C32 a_n1665_109# a_n1949_109# 0.06fF
C33 a_n1089_109# a_n1089_527# 0.01fF
C34 a_n33_n309# a_n33_109# 0.01fF
C35 a_831_527# a_831_109# 0.01fF
C36 a_1791_n309# a_1695_n309# 0.29fF
C37 a_63_109# a_351_109# 0.06fF
C38 a_1215_n309# a_1407_n309# 0.11fF
C39 a_447_527# a_447_109# 0.01fF
C40 a_n801_527# a_n1185_527# 0.05fF
C41 a_1119_n309# a_1119_109# 0.01fF
C42 a_n225_n309# a_n225_109# 0.01fF
C43 a_1503_n309# a_1119_n309# 0.05fF
C44 a_n993_109# a_n1377_109# 0.05fF
C45 a_159_109# a_n129_109# 0.06fF
C46 a_n705_109# a_n897_109# 0.11fF
C47 a_n225_527# a_n225_109# 0.01fF
C48 a_n801_n309# a_n1089_n309# 0.06fF
C49 a_n225_n727# a_n417_n727# 0.11fF
C50 a_735_109# a_735_n309# 0.01fF
C51 a_n993_109# a_n1089_109# 0.29fF
C52 a_1887_n727# a_1503_n727# 0.05fF
C53 a_n129_n309# a_255_n309# 0.05fF
C54 a_n1185_527# a_n993_527# 0.11fF
C55 a_1599_109# a_1887_109# 0.06fF
C56 a_n321_109# a_n417_109# 0.29fF
C57 a_1407_527# a_1023_527# 0.05fF
C58 a_1887_n309# a_1887_n727# 0.01fF
C59 a_159_527# a_351_527# 0.11fF
C60 a_735_527# a_351_527# 0.05fF
C61 a_63_n309# a_n321_n309# 0.05fF
C62 a_n609_109# a_n513_109# 0.29fF
C63 a_447_527# a_63_527# 0.05fF
C64 a_1215_n309# a_1119_n309# 0.29fF
C65 a_1503_n309# a_1695_n309# 0.11fF
C66 a_831_n309# a_735_n309# 0.29fF
C67 a_n1569_527# a_n1377_527# 0.11fF
C68 a_255_n727# a_159_n727# 0.29fF
C69 a_1119_n727# a_1023_n727# 0.29fF
C70 a_543_527# a_927_527# 0.05fF
C71 a_639_n309# a_351_n309# 0.06fF
C72 a_n33_n727# a_n417_n727# 0.05fF
C73 a_n1281_n727# a_n1665_n727# 0.05fF
C74 a_447_n727# a_351_n727# 0.29fF
C75 a_1695_109# a_1695_n309# 0.01fF
C76 a_1407_n309# a_1023_n309# 0.05fF
C77 a_543_109# a_255_109# 0.06fF
C78 a_1119_n727# a_1311_n727# 0.11fF
C79 a_447_109# a_255_109# 0.11fF
C80 a_1215_n309# a_927_n309# 0.06fF
C81 a_n1089_n727# a_n1089_n309# 0.01fF
C82 a_n897_109# a_n897_n309# 0.01fF
C83 a_n609_n309# a_n225_n309# 0.05fF
C84 a_255_n309# a_255_109# 0.01fF
C85 a_447_n727# a_63_n727# 0.05fF
C86 a_1503_527# a_1215_527# 0.06fF
C87 a_n513_n727# a_n417_n727# 0.29fF
C88 a_159_527# a_159_109# 0.01fF
C89 a_n1089_109# a_n1377_109# 0.06fF
C90 a_n513_527# a_n321_527# 0.11fF
C91 a_n1185_109# a_n993_109# 0.11fF
C92 a_831_527# a_1215_527# 0.05fF
C93 a_n897_n309# a_n1185_n309# 0.06fF
C94 a_n129_n309# a_n129_n727# 0.01fF
C95 a_n1569_527# a_n1185_527# 0.05fF
C96 a_1791_109# a_1791_527# 0.01fF
C97 a_n1185_n727# a_n1089_n727# 0.29fF
C98 a_n897_527# a_n1089_527# 0.11fF
C99 a_n1857_n727# a_n1761_n727# 0.29fF
C100 a_n993_n309# a_n705_n309# 0.06fF
C101 a_n1665_109# a_n1377_109# 0.06fF
C102 a_543_527# a_159_527# 0.05fF
C103 a_927_n727# a_1215_n727# 0.06fF
C104 a_543_527# a_735_527# 0.11fF
C105 a_639_n309# a_255_n309# 0.05fF
C106 a_n321_109# a_n33_109# 0.06fF
C107 a_n225_527# a_n33_527# 0.11fF
C108 a_1023_n309# a_1119_n309# 0.29fF
C109 a_n1665_527# a_n1949_527# 0.06fF
C110 a_1407_527# a_1407_109# 0.01fF
C111 a_1311_n309# a_1311_109# 0.01fF
C112 a_n321_527# a_n609_527# 0.06fF
C113 a_n1377_n309# a_n993_n309# 0.05fF
C114 a_1407_n309# a_1119_n309# 0.06fF
C115 a_831_527# a_639_527# 0.11fF
C116 a_1119_527# a_1119_109# 0.01fF
C117 a_n321_527# a_n321_109# 0.01fF
C118 a_n33_n309# a_n225_n309# 0.11fF
C119 a_543_n309# a_831_n309# 0.06fF
C120 a_n1281_n309# a_n993_n309# 0.06fF
C121 a_n1949_n727# a_n1569_n727# 0.05fF
C122 a_447_n727# a_543_n727# 0.29fF
C123 a_1023_n309# a_927_n309# 0.29fF
C124 a_n225_n727# a_63_n727# 0.06fF
C125 a_n1569_109# a_n1569_n309# 0.01fF
C126 a_n609_n309# a_n993_n309# 0.05fF
C127 a_n513_n309# a_n897_n309# 0.05fF
C128 a_639_n309# a_1023_n309# 0.05fF
C129 a_n1281_527# a_n1665_527# 0.05fF
C130 a_n1185_109# a_n1377_109# 0.11fF
C131 a_n609_109# a_n801_109# 0.11fF
C132 a_351_n309# a_63_n309# 0.06fF
C133 a_n33_n727# a_351_n727# 0.05fF
C134 a_n1569_n727# a_n1665_n727# 0.29fF
C135 a_n801_527# a_n1089_527# 0.06fF
C136 a_n1569_109# a_n1281_109# 0.06fF
C137 a_n1185_109# a_n1089_109# 0.29fF
C138 a_639_527# a_255_527# 0.05fF
C139 a_n1185_n727# a_n1377_n727# 0.11fF
C140 a_n513_527# a_n609_527# 0.29fF
C141 a_255_n727# a_255_n309# 0.01fF
C142 a_1407_n309# a_1695_n309# 0.06fF
C143 a_n1089_n727# a_n1377_n727# 0.06fF
C144 a_n1473_n727# a_n1761_n727# 0.06fF
C145 a_n33_n727# a_63_n727# 0.29fF
C146 a_255_527# a_n33_527# 0.06fF
C147 a_351_109# a_n33_109# 0.05fF
C148 a_1407_527# a_1215_527# 0.11fF
C149 a_1599_n727# a_1503_n727# 0.29fF
C150 a_n321_n727# a_n417_n727# 0.29fF
C151 a_735_109# a_1119_109# 0.05fF
C152 a_n417_527# a_n417_109# 0.01fF
C153 a_639_n309# a_639_n727# 0.01fF
C154 a_n1473_527# a_n1281_527# 0.11fF
C155 a_n513_n309# a_n321_n309# 0.11fF
C156 a_n1857_n309# a_n1569_n309# 0.06fF
C157 a_n1089_527# a_n993_527# 0.29fF
C158 a_n1761_109# a_n1761_n309# 0.01fF
C159 a_n321_527# a_n225_527# 0.29fF
C160 a_n1473_109# a_n1377_109# 0.29fF
C161 a_n993_109# a_n993_n309# 0.01fF
C162 a_1887_527# a_1887_109# 0.01fF
C163 a_n129_n309# a_n129_109# 0.01fF
C164 a_n1473_109# a_n1089_109# 0.05fF
C165 a_927_n727# a_1119_n727# 0.11fF
C166 a_n993_n727# a_n609_n727# 0.05fF
C167 a_n417_527# a_n33_527# 0.05fF
C168 a_1119_n309# a_927_n309# 0.11fF
C169 a_255_n309# a_63_n309# 0.11fF
C170 a_n1665_527# a_n1377_527# 0.06fF
C171 a_1695_n727# a_1503_n727# 0.11fF
C172 a_n609_109# a_n897_109# 0.06fF
C173 a_n1473_109# a_n1665_109# 0.11fF
C174 a_n993_109# a_n993_527# 0.01fF
C175 a_n1949_527# a_n1761_527# 0.11fF
C176 a_1407_n309# a_1407_n727# 0.01fF
C177 a_n801_n309# a_n801_109# 0.01fF
C178 a_n513_527# a_n897_527# 0.05fF
C179 a_1119_n727# a_1215_n727# 0.29fF
C180 a_n513_527# a_n225_527# 0.06fF
C181 a_n993_n727# a_n897_n727# 0.29fF
C182 a_n417_n309# a_n321_n309# 0.29fF
C183 a_n1473_n309# a_n1089_n309# 0.05fF
C184 a_255_n727# a_n129_n727# 0.05fF
C185 a_1311_527# a_927_527# 0.05fF
C186 a_255_n727# a_639_n727# 0.05fF
C187 a_639_n727# a_735_n727# 0.29fF
C188 a_639_n309# a_927_n309# 0.06fF
C189 a_1215_n309# a_831_n309# 0.05fF
C190 a_735_109# a_543_109# 0.11fF
C191 a_1599_n727# a_1599_n309# 0.01fF
C192 a_735_109# a_447_109# 0.06fF
C193 a_735_527# a_447_527# 0.06fF
C194 a_159_527# a_447_527# 0.06fF
C195 a_1311_n727# a_1503_n727# 0.11fF
C196 a_159_527# a_63_527# 0.29fF
C197 a_255_109# a_n129_109# 0.05fF
C198 a_n1473_527# a_n1377_527# 0.29fF
C199 a_n609_n727# a_n801_n727# 0.11fF
C200 a_n705_n727# a_n417_n727# 0.06fF
C201 a_1215_527# a_1599_527# 0.05fF
C202 a_n129_n309# a_63_n309# 0.11fF
C203 a_n897_527# a_n609_527# 0.06fF
C204 a_n225_527# a_n609_527# 0.05fF
C205 a_n1185_109# a_n1473_109# 0.06fF
C206 a_1311_n309# a_1311_n727# 0.01fF
C207 a_447_n727# a_159_n727# 0.06fF
C208 a_n705_109# a_n705_n309# 0.01fF
C209 a_n513_109# a_n129_109# 0.05fF
C210 a_n897_n727# a_n801_n727# 0.29fF
C211 a_n321_527# a_n417_527# 0.29fF
C212 a_1119_527# a_1311_527# 0.11fF
C213 a_n1473_n727# a_n1281_n727# 0.11fF
C214 a_639_n727# a_831_n727# 0.11fF
C215 a_n513_527# a_n801_527# 0.06fF
C216 a_n321_n727# a_63_n727# 0.05fF
C217 a_n1473_527# a_n1185_527# 0.06fF
C218 a_159_n309# a_543_n309# 0.05fF
C219 a_n1569_n309# a_n1473_n309# 0.29fF
C220 a_n1569_n309# a_n1949_n309# 0.05fF
C221 a_159_n309# a_159_109# 0.01fF
C222 a_n1949_n727# a_n1665_n727# 0.06fF
C223 a_n1761_109# a_n1949_109# 0.11fF
C224 a_n1857_n309# a_n1473_n309# 0.05fF
C225 a_n705_109# a_n417_109# 0.06fF
C226 a_n1857_n309# a_n1949_n309# 0.29fF
C227 a_1023_n309# a_831_n309# 0.11fF
C228 a_n1857_n727# a_n1569_n727# 0.06fF
C229 a_n801_n309# a_n1185_n309# 0.05fF
C230 a_n801_527# a_n609_527# 0.11fF
C231 a_n513_527# a_n417_527# 0.29fF
C232 a_1311_109# a_1503_109# 0.11fF
C233 a_159_n309# a_159_n727# 0.01fF
C234 a_1887_n309# a_1887_109# 0.01fF
C235 a_n897_n309# a_n705_n309# 0.11fF
C236 a_n1761_527# a_n1377_527# 0.05fF
C237 a_n1089_n309# a_n1185_n309# 0.29fF
C238 a_n225_n727# a_159_n727# 0.05fF
C239 a_1311_109# a_1119_109# 0.11fF
C240 a_n1949_109# a_n1857_109# 0.29fF
C241 a_n513_109# a_n801_109# 0.06fF
C242 a_1791_n727# a_1503_n727# 0.06fF
C243 a_n609_527# a_n993_527# 0.05fF
C244 a_63_109# a_159_109# 0.29fF
C245 a_n1185_n727# a_n993_n727# 0.11fF
C246 a_n801_n309# a_n801_n727# 0.01fF
C247 a_n993_n727# a_n1089_n727# 0.29fF
C248 a_n417_527# a_n609_527# 0.11fF
C249 a_n1185_n727# a_n1185_n309# 0.01fF
C250 a_543_109# a_639_109# 0.29fF
C251 a_n1281_n309# a_n897_n309# 0.05fF
C252 a_n225_n727# a_n609_n727# 0.05fF
C253 a_n705_n309# a_n321_n309# 0.05fF
C254 a_n33_n727# a_159_n727# 0.11fF
C255 a_447_109# a_639_109# 0.11fF
C256 a_1311_109# a_1695_109# 0.05fF
C257 a_n993_109# a_n705_109# 0.06fF
C258 a_1215_109# a_1503_109# 0.06fF
C259 a_n801_n309# a_n513_n309# 0.06fF
C260 a_n609_n309# a_n897_n309# 0.06fF
C261 a_1119_n309# a_831_n309# 0.06fF
C262 a_159_109# a_n225_109# 0.05fF
C263 a_1215_109# a_1119_109# 0.29fF
C264 a_n801_527# a_n897_527# 0.29fF
C265 a_831_109# a_1119_109# 0.06fF
C266 a_159_n309# a_351_n309# 0.11fF
C267 a_n1473_n727# a_n1569_n727# 0.29fF
C268 a_1119_527# a_927_527# 0.11fF
C269 a_n897_109# a_n1281_109# 0.05fF
C270 a_1023_109# a_1119_109# 0.29fF
C271 a_n1185_n727# a_n801_n727# 0.05fF
C272 a_63_527# a_n129_527# 0.11fF
C273 a_1887_527# a_1503_527# 0.05fF
C274 a_735_527# a_927_527# 0.11fF
C275 a_831_n309# a_927_n309# 0.29fF
C276 a_n1569_n309# a_n1185_n309# 0.05fF
C277 a_n1089_n727# a_n801_n727# 0.06fF
C278 a_1791_109# a_1791_n309# 0.01fF
C279 a_n609_n309# a_n321_n309# 0.06fF
C280 a_n513_n309# a_n129_n309# 0.05fF
C281 a_1503_109# a_1407_109# 0.29fF
C282 a_735_n727# a_831_n727# 0.29fF
C283 a_1503_527# a_1791_527# 0.06fF
C284 a_639_n309# a_831_n309# 0.11fF
C285 a_n897_527# a_n993_527# 0.29fF
C286 a_n897_109# a_n513_109# 0.05fF
C287 a_1503_n727# a_1215_n727# 0.06fF
C288 a_1599_109# a_1599_527# 0.01fF
C289 a_639_527# a_351_527# 0.06fF
C290 a_n801_n309# a_n417_n309# 0.05fF
C291 a_n993_n727# a_n1377_n727# 0.05fF
C292 a_1407_109# a_1119_109# 0.06fF
C293 a_n417_527# a_n225_527# 0.11fF
C294 a_1215_n309# a_1215_109# 0.01fF
C295 a_351_527# a_n33_527# 0.05fF
C296 a_n513_n727# a_n609_n727# 0.29fF
C297 a_n321_n727# a_n321_n309# 0.01fF
C298 a_n1761_109# a_n1377_109# 0.05fF
C299 a_n1281_527# a_n1281_109# 0.01fF
C300 a_n705_109# a_n1089_109# 0.05fF
C301 a_1791_109# a_1503_109# 0.06fF
C302 a_159_n309# a_255_n309# 0.29fF
C303 a_735_527# a_1119_527# 0.05fF
C304 a_543_109# a_831_109# 0.06fF
C305 a_1695_109# a_1407_109# 0.06fF
C306 a_n609_109# a_n225_109# 0.05fF
C307 a_927_n727# a_543_n727# 0.05fF
C308 a_831_109# a_447_109# 0.05fF
C309 a_1887_527# a_1791_527# 0.29fF
C310 a_n513_n727# a_n897_n727# 0.05fF
C311 a_1407_527# a_1503_527# 0.29fF
C312 a_n129_n309# a_n417_n309# 0.06fF
C313 a_n1473_527# a_n1089_527# 0.05fF
C314 a_639_n727# a_447_n727# 0.11fF
C315 a_1599_109# a_1599_n309# 0.01fF
C316 a_n1665_109# a_n1761_109# 0.29fF
C317 a_n1857_n727# a_n1949_n727# 0.29fF
C318 a_n801_527# a_n993_527# 0.11fF
C319 a_n33_n309# a_n321_n309# 0.06fF
C320 a_63_109# a_447_109# 0.05fF
C321 a_639_109# a_255_109# 0.05fF
C322 a_n801_527# a_n417_527# 0.05fF
C323 a_1791_109# a_1695_109# 0.29fF
C324 a_n1857_n727# a_n1665_n727# 0.11fF
C325 a_n513_n309# a_n513_109# 0.01fF
C326 a_543_527# a_639_527# 0.29fF
C327 a_1311_527# a_1023_527# 0.06fF
C328 a_1311_109# a_1311_527# 0.01fF
C329 a_n897_n727# a_n1281_n727# 0.05fF
C330 a_735_527# a_735_109# 0.01fF
C331 a_159_n309# a_n129_n309# 0.06fF
C332 a_n1665_109# a_n1857_109# 0.11fF
C333 a_n609_n309# a_n609_n727# 0.01fF
C334 a_n705_109# a_n321_109# 0.05fF
C335 a_1119_n727# a_1503_n727# 0.05fF
C336 a_1407_527# a_1791_527# 0.05fF
C337 a_639_n309# a_639_109# 0.01fF
C338 a_1023_n309# a_1023_109# 0.01fF
C339 a_n321_n727# a_n609_n727# 0.06fF
C340 a_63_109# a_63_527# 0.01fF
C341 a_n609_109# a_n417_109# 0.11fF
C342 a_831_n727# a_831_n309# 0.01fF
C343 a_n225_n727# a_n129_n727# 0.29fF
C344 a_n609_109# a_n609_n309# 0.01fF
C345 a_1695_527# a_1503_527# 0.11fF
C346 a_n897_109# a_n801_109# 0.29fF
C347 a_n1569_n309# a_n1665_n309# 0.29fF
C348 a_159_109# a_n33_109# 0.11fF
C349 a_n1473_n309# a_n1185_n309# 0.06fF
C350 a_n1857_n309# a_n1665_n309# 0.11fF
C351 a_n129_109# a_n129_527# 0.01fF
C352 a_1791_n727# a_1791_n309# 0.01fF
C353 a_1503_527# a_1599_527# 0.29fF
C354 a_1503_109# a_1887_109# 0.05fF
C355 a_n33_n727# a_n129_n727# 0.29fF
C356 a_n1473_109# a_n1761_109# 0.06fF
C357 a_n1569_n309# a_n1761_n309# 0.11fF
C358 a_1407_n309# a_1407_109# 0.01fF
C359 a_n801_n309# a_n705_n309# 0.29fF
C360 a_n1473_n727# a_n1665_n727# 0.11fF
C361 a_n1857_n309# a_n1761_n309# 0.29fF
C362 a_n1665_527# a_n1665_109# 0.01fF
C363 a_1695_527# a_1887_527# 0.11fF
C364 a_n1377_n727# a_n1761_n727# 0.05fF
C365 a_n1089_n309# a_n705_n309# 0.05fF
C366 a_n609_109# a_n993_109# 0.05fF
C367 a_1695_527# a_1791_527# 0.29fF
C368 a_n513_n727# a_n129_n727# 0.05fF
C369 a_n1473_109# a_n1857_109# 0.05fF
C370 a_735_n727# a_447_n727# 0.06fF
C371 a_255_n727# a_447_n727# 0.11fF
C372 a_1887_527# a_1599_527# 0.06fF
C373 a_63_109# a_255_109# 0.11fF
C374 a_351_n309# a_n33_n309# 0.05fF
C375 a_1023_n309# a_1023_n727# 0.01fF
C376 a_1695_109# a_1887_109# 0.11fF
C377 a_1791_527# a_1599_527# 0.11fF
C378 a_n321_109# a_n321_n309# 0.01fF
C379 a_n1089_n309# a_n1377_n309# 0.06fF
C380 a_n801_n309# a_n609_n309# 0.11fF
C381 a_n1857_527# a_n1569_527# 0.06fF
C382 a_927_527# a_1023_527# 0.29fF
C383 a_n705_n727# a_n609_n727# 0.29fF
C384 a_447_n309# a_735_n309# 0.06fF
C385 a_n1281_n309# a_n1089_n309# 0.11fF
C386 a_159_527# a_n129_527# 0.06fF
C387 a_n1185_n727# a_n1281_n727# 0.29fF
C388 a_n1089_n727# a_n1281_n727# 0.11fF
C389 a_639_n727# a_1023_n727# 0.05fF
C390 a_1407_527# a_1695_527# 0.06fF
C391 a_1599_109# a_1503_109# 0.29fF
C392 a_n705_n727# a_n897_n727# 0.11fF
C393 a_639_527# a_447_527# 0.11fF
C394 a_447_n727# a_831_n727# 0.05fF
C395 a_1311_527# a_1215_527# 0.29fF
C396 a_n225_n309# a_n321_n309# 0.29fF
C397 a_1407_527# a_1599_527# 0.11fF
C398 a_n33_527# a_63_527# 0.29fF
C399 a_n513_109# a_n225_109# 0.06fF
C400 a_n1569_109# a_n1949_109# 0.05fF
C401 a_255_n309# a_n33_n309# 0.06fF
C402 a_1119_527# a_1023_527# 0.29fF
C403 a_351_527# a_351_109# 0.01fF
C404 a_735_109# a_639_109# 0.29fF
C405 a_735_527# a_1023_527# 0.06fF
C406 a_n1949_n309# a_n1665_n309# 0.06fF
C407 a_63_109# a_n129_109# 0.11fF
C408 a_n1473_n309# a_n1665_n309# 0.11fF
C409 a_n993_n727# a_n801_n727# 0.11fF
C410 a_1695_109# a_1599_109# 0.29fF
C411 a_n1569_n309# a_n1377_n309# 0.11fF
C412 a_n321_n727# a_n129_n727# 0.11fF
C413 a_n897_n309# a_n993_n309# 0.29fF
C414 a_n1473_527# a_n1473_109# 0.01fF
C415 a_n33_n727# a_255_n727# 0.06fF
C416 a_1695_n727# a_1695_n309# 0.01fF
C417 a_n1281_n309# a_n1569_n309# 0.06fF
C418 a_n1377_n727# a_n1281_n727# 0.29fF
C419 a_n1949_n309# a_n1761_n309# 0.11fF
C420 a_n1473_n309# a_n1761_n309# 0.06fF
C421 a_159_n309# a_63_n309# 0.29fF
C422 a_63_n727# a_351_n727# 0.06fF
C423 a_n129_109# a_n225_109# 0.29fF
C424 a_n1281_n309# a_n1281_109# 0.01fF
C425 a_1599_n727# a_1407_n727# 0.11fF
C426 a_1215_n309# a_1215_n727# 0.01fF
C427 a_n129_n309# a_n33_n309# 0.29fF
C428 a_n1377_n727# a_n1377_n309# 0.01fF
C429 a_351_109# a_159_109# 0.11fF
C430 a_543_n309# a_447_n309# 0.29fF
C431 a_n609_109# a_n609_527# 0.01fF
C432 a_351_527# a_255_527# 0.29fF
C433 a_1695_527# a_1599_527# 0.29fF
C434 a_n609_109# a_n321_109# 0.06fF
C435 a_n513_109# a_n417_109# 0.29fF
C436 a_n1857_527# a_n1857_109# 0.01fF
C437 a_n1185_n727# a_n1569_n727# 0.05fF
C438 a_n1857_n727# a_n1473_n727# 0.05fF
C439 a_n321_527# a_63_527# 0.05fF
C440 a_63_109# a_63_n309# 0.01fF
C441 a_927_109# a_1119_109# 0.11fF
C442 a_1695_n727# a_1407_n727# 0.06fF
C443 a_n1281_527# a_n1377_527# 0.29fF
C444 a_n1089_109# a_n1089_n309# 0.01fF
C445 a_735_109# a_831_109# 0.29fF
C446 a_543_527# a_831_527# 0.06fF
C447 a_735_n727# a_1023_n727# 0.06fF
C448 a_927_527# a_1215_527# 0.06fF
C449 a_351_n727# a_543_n727# 0.11fF
C450 a_1407_n727# a_1023_n727# 0.05fF
C451 a_n993_109# a_n1281_109# 0.06fF
C452 a_1503_527# a_1503_109# 0.01fF
C453 a_735_109# a_1023_109# 0.06fF
C454 a_n705_n727# a_n1089_n727# 0.05fF
C455 a_n417_109# a_n129_109# 0.06fF
C456 a_n1569_n309# a_n1569_n727# 0.01fF
C457 a_831_109# a_831_n309# 0.01fF
C458 a_1887_n309# a_1599_n309# 0.06fF
C459 a_1311_n727# a_1407_n727# 0.29fF
C460 a_255_109# a_n33_109# 0.06fF
C461 a_n1569_109# a_n1377_109# 0.11fF
C462 a_927_n727# a_639_n727# 0.06fF
C463 a_351_n309# a_351_109# 0.01fF
C464 a_1311_n309# a_1599_n309# 0.06fF
C465 a_n1857_527# a_n1665_527# 0.11fF
C466 a_447_n309# a_351_n309# 0.29fF
C467 a_543_527# a_255_527# 0.06fF
C468 a_n705_527# a_n1089_527# 0.05fF
C469 a_n1281_527# a_n1185_527# 0.29fF
C470 a_n1377_n727# a_n1569_n727# 0.11fF
C471 a_639_527# a_927_527# 0.06fF
C472 a_1119_527# a_1215_527# 0.29fF
C473 a_n513_n309# a_n417_n309# 0.29fF
C474 a_831_n727# a_1023_n727# 0.11fF
C475 a_543_109# a_927_109# 0.05fF
C476 a_n1473_n309# a_n1377_n309# 0.29fF
C477 a_n1569_109# a_n1665_109# 0.29fF
C478 a_n609_n727# a_n417_n727# 0.11fF
C479 a_n1949_n309# a_n1949_109# 0.01fF
C480 a_n1281_n309# a_n1473_n309# 0.11fF
C481 a_n1665_527# a_n1569_527# 0.29fF
C482 a_n1473_527# a_n1857_527# 0.05fF
C483 a_n1281_109# a_n1377_109# 0.29fF
C484 a_543_109# a_351_109# 0.11fF
C485 a_n1089_109# a_n1281_109# 0.11fF
C486 a_351_109# a_447_109# 0.29fF
C487 a_n801_109# a_n417_109# 0.05fF
C488 a_n1761_109# a_n1857_109# 0.29fF
C489 a_447_n309# a_447_109# 0.01fF
C490 a_927_n727# a_927_n309# 0.01fF
C491 a_255_n309# a_447_n309# 0.11fF
C492 a_n129_109# a_n33_109# 0.29fF
C493 a_n1473_527# a_n1569_527# 0.29fF
C494 a_735_527# a_639_527# 0.29fF
C495 a_n1665_109# a_n1281_109# 0.05fF
C496 a_n1569_109# a_n1185_109# 0.05fF
C497 a_159_527# a_n33_527# 0.11fF
C498 a_n1185_527# a_n1377_527# 0.11fF
C499 a_n513_527# a_n513_109# 0.01fF
C500 a_1599_n727# a_1887_n727# 0.06fF
C501 a_1791_n727# a_1407_n727# 0.05fF
C502 a_n225_527# a_63_527# 0.06fF
C503 a_831_109# a_639_109# 0.11fF
C504 a_n129_n309# a_n225_n309# 0.29fF
C505 a_n993_n727# a_n1281_n727# 0.06fF
C506 a_n705_527# a_n321_527# 0.05fF
C507 a_639_109# a_1023_109# 0.05fF
C508 a_159_n727# a_351_n727# 0.11fF
C509 a_n993_109# a_n801_109# 0.11fF
C510 a_n513_n727# a_n801_n727# 0.06fF
C511 a_63_n309# a_n33_n309# 0.29fF
C512 a_831_527# a_447_527# 0.05fF
C513 a_n1569_109# a_n1473_109# 0.29fF
C514 a_n1857_527# a_n1761_527# 0.29fF
C515 a_n1949_527# a_n1949_109# 0.01fF
C516 a_n1185_109# a_n1281_109# 0.29fF
C517 a_159_n727# a_63_n727# 0.29fF
C518 a_927_n727# a_735_n727# 0.11fF
C519 a_1887_n309# a_1791_n309# 0.29fF
C520 a_n1185_n309# a_n1377_n309# 0.11fF
C521 a_n513_n309# a_n513_n727# 0.01fF
C522 a_n801_n309# a_n993_n309# 0.11fF
C523 a_1311_109# a_1215_109# 0.29fF
C524 a_n321_109# a_n513_109# 0.11fF
C525 a_1695_n727# a_1887_n727# 0.11fF
C526 a_n1761_n309# a_n1665_n309# 0.29fF
C527 a_n1281_n309# a_n1185_n309# 0.29fF
C528 a_n705_527# a_n513_527# 0.11fF
C529 a_1311_109# a_1023_109# 0.06fF
C530 a_n1089_n309# a_n993_n309# 0.29fF
C531 a_1023_527# a_1023_109# 0.01fF
C532 a_n1761_n309# a_n1761_n727# 0.01fF
C533 a_1311_527# a_1503_527# 0.11fF
C534 a_n1569_527# a_n1761_527# 0.11fF
C535 a_447_527# a_255_527# 0.11fF
C536 a_255_527# a_63_527# 0.11fF
C537 a_1119_n727# a_1119_n309# 0.01fF
C538 a_n513_n309# a_n705_n309# 0.11fF
C539 a_n1473_109# a_n1281_109# 0.11fF
C540 a_1407_n727# a_1215_n727# 0.11fF
C541 a_351_109# a_255_109# 0.29fF
C542 a_351_n309# a_351_n727# 0.01fF
C543 a_1503_n309# a_1503_n727# 0.01fF
C544 a_543_n309# a_543_n727# 0.01fF
C545 a_927_109# a_927_n309# 0.01fF
C546 a_1311_109# a_1407_109# 0.29fF
C547 a_n321_109# a_n129_109# 0.11fF
C548 a_1887_n309# a_1503_n309# 0.05fF
C549 a_927_n727# a_831_n727# 0.29fF
C550 a_n705_527# a_n609_527# 0.29fF
C551 a_831_109# a_1215_109# 0.05fF
C552 a_n1281_527# a_n1089_527# 0.11fF
C553 a_n993_109# a_n897_109# 0.29fF
C554 a_n801_109# a_n1089_109# 0.06fF
C555 a_543_n309# a_735_n309# 0.11fF
C556 a_1791_n309# a_1599_n309# 0.11fF
C557 a_1311_n309# a_1503_n309# 0.11fF
C558 a_n1377_n727# a_n1665_n727# 0.06fF
C559 a_n129_n727# a_n417_n727# 0.06fF
C560 a_159_n727# a_543_n727# 0.05fF
C561 a_1695_527# a_1695_109# 0.01fF
C562 a_1215_109# a_1023_109# 0.11fF
C563 a_n33_n727# a_n225_n727# 0.11fF
C564 a_831_109# a_1023_109# 0.11fF
C565 a_n513_n309# a_n609_n309# 0.29fF
C566 a_639_n309# a_447_n309# 0.11fF
C567 a_831_n727# a_1215_n727# 0.05fF
C568 a_n417_n309# a_n705_n309# 0.06fF
C569 a_1215_109# a_1407_109# 0.11fF
C570 a_1215_n309# a_1311_n309# 0.29fF
C571 a_n225_n727# a_n513_n727# 0.06fF
C572 a_n609_109# a_n705_109# 0.29fF
C573 a_255_527# a_255_109# 0.01fF
C574 a_927_527# a_927_109# 0.01fF
C575 a_n1761_109# a_n1761_527# 0.01fF
C576 a_1023_109# a_1407_109# 0.05fF
C577 a_1023_527# a_1215_527# 0.11fF
C578 a_639_527# a_639_109# 0.01fF
C579 a_n33_527# a_n129_527# 0.29fF
C580 a_1503_n309# a_1599_n309# 0.29fF
C581 a_n705_n727# a_n993_n727# 0.06fF
C582 a_n705_527# a_n897_527# 0.11fF
C583 a_n1473_527# a_n1665_527# 0.11fF
C584 a_1407_527# a_1311_527# 0.29fF
C585 a_n417_n309# a_n417_109# 0.01fF
C586 a_n1089_527# a_n1377_527# 0.06fF
C587 a_n1185_109# a_n801_109# 0.05fF
C588 a_1119_n727# a_735_n727# 0.05fF
C589 a_n897_109# a_n1089_109# 0.11fF
C590 a_n417_n309# a_n609_n309# 0.11fF
C591 a_n1665_n309# a_n1377_n309# 0.06fF
C592 a_1119_n727# a_1407_n727# 0.06fF
C593 a_63_109# a_n225_109# 0.06fF
C594 a_1791_n727# a_1887_n727# 0.29fF
C595 a_n1281_n309# a_n1665_n309# 0.05fF
C596 a_543_527# a_351_527# 0.11fF
C597 a_351_n309# a_735_n309# 0.05fF
C598 a_1215_n309# a_1599_n309# 0.05fF
C599 a_n1949_n727# a_n1949_n309# 0.01fF
C600 a_639_527# a_1023_527# 0.05fF
C601 a_831_527# a_927_527# 0.29fF
C602 a_n1761_n309# a_n1377_n309# 0.05fF
C603 a_1215_109# a_1215_527# 0.01fF
C604 a_n1473_109# a_n1473_n309# 0.01fF
C605 a_63_n309# a_n225_n309# 0.06fF
C606 a_n897_n309# a_n897_n727# 0.01fF
C607 a_n1569_109# a_n1569_527# 0.01fF
C608 a_1599_n727# a_1695_n727# 0.29fF
C609 a_1791_109# a_1407_109# 0.05fF
C610 a_n705_n727# a_n801_n727# 0.29fF
C611 a_n1185_527# a_n1089_527# 0.29fF
C612 a_1311_n309# a_1023_n309# 0.06fF
C613 a_639_n727# a_351_n727# 0.06fF
C614 a_1119_n727# a_831_n727# 0.06fF
C615 a_n705_527# a_n801_527# 0.29fF
C616 a_159_527# a_n225_527# 0.05fF
C617 a_1119_527# a_1503_527# 0.05fF
C618 a_447_n309# a_63_n309# 0.05fF
C619 a_n129_n727# a_63_n727# 0.11fF
C620 a_n321_527# a_n129_527# 0.11fF
C621 a_1311_n309# a_1407_n309# 0.29fF
C622 a_n417_n309# a_n33_n309# 0.05fF
C623 a_1695_527# a_1311_527# 0.05fF
C624 a_n321_n727# a_n225_n727# 0.29fF
C625 a_831_527# a_1119_527# 0.06fF
C626 a_n1185_109# a_n897_109# 0.06fF
C627 a_1599_n727# a_1311_n727# 0.06fF
C628 a_735_109# a_927_109# 0.11fF
C629 a_n1665_527# a_n1761_527# 0.29fF
C630 a_n1857_n727# a_n1857_n309# 0.01fF
C631 a_n705_527# a_n993_527# 0.06fF
C632 a_831_527# a_735_527# 0.29fF
C633 a_1311_527# a_1599_527# 0.06fF
C634 a_n705_527# a_n417_527# 0.06fF
C635 a_n1185_109# a_n1185_n309# 0.01fF
C636 a_735_109# a_351_109# 0.05fF
C637 a_n33_n727# a_n321_n727# 0.06fF
C638 a_n1377_109# a_n1377_527# 0.01fF
C639 a_n1185_n727# a_n1473_n727# 0.06fF
C640 a_159_n309# a_n33_n309# 0.11fF
C641 a_n1089_n727# a_n1473_n727# 0.05fF
C642 a_n1569_n727# a_n1761_n727# 0.11fF
C643 a_n417_109# a_n225_109# 0.11fF
C644 a_n513_527# a_n129_527# 0.05fF
C645 a_n801_527# a_n801_109# 0.01fF
C646 a_n1473_527# a_n1761_527# 0.06fF
C647 a_543_n309# a_351_n309# 0.11fF
C648 a_1311_n309# a_1119_n309# 0.11fF
C649 a_n801_n309# a_n897_n309# 0.29fF
C650 a_1407_n309# a_1599_n309# 0.11fF
C651 a_1023_n309# a_735_n309# 0.06fF
C652 a_159_527# a_255_527# 0.29fF
C653 a_n1569_109# a_n1761_109# 0.11fF
C654 a_1311_n727# a_1695_n727# 0.05fF
C655 a_1503_n309# a_1791_n309# 0.06fF
C656 a_n897_109# a_n897_527# 0.01fF
C657 a_447_n309# a_831_n309# 0.05fF
C658 a_n1089_n309# a_n897_n309# 0.11fF
C659 a_1311_n727# a_1023_n727# 0.06fF
C660 a_n321_n727# a_n513_n727# 0.11fF
C661 a_639_n727# a_543_n727# 0.29fF
C662 a_1887_n309# a_1695_n309# 0.11fF
C663 a_n609_n309# a_n705_n309# 0.29fF
C664 a_1311_n309# a_927_n309# 0.05fF
C665 a_n1281_n309# a_n1281_n727# 0.01fF
C666 a_1311_109# a_1599_109# 0.06fF
C667 a_n33_n727# a_n33_n309# 0.01fF
C668 a_1503_109# a_1119_109# 0.05fF
C669 a_n1569_109# a_n1857_109# 0.06fF
C670 a_1311_n309# a_1695_n309# 0.05fF
C671 a_1503_n309# a_1503_109# 0.01fF
C672 a_n1281_n309# a_n1377_n309# 0.29fF
C673 a_1407_527# a_1119_527# 0.06fF
C674 a_351_527# a_447_527# 0.29fF
C675 a_n1281_527# a_n897_527# 0.05fF
C676 a_543_n309# a_543_109# 0.01fF
C677 a_63_109# a_n33_109# 0.29fF
C678 a_n609_n727# a_n897_n727# 0.06fF
C679 a_351_527# a_63_527# 0.06fF
C680 a_543_109# a_159_109# 0.05fF
C681 a_1599_n727# a_1791_n727# 0.11fF
C682 a_447_109# a_159_109# 0.06fF
C683 a_543_n309# a_255_n309# 0.06fF
C684 a_n1665_109# a_n1665_n309# 0.01fF
C685 a_n705_109# a_n513_109# 0.11fF
C686 a_n1473_n727# a_n1377_n727# 0.29fF
C687 a_1695_109# a_1503_109# 0.11fF
C688 a_255_n727# a_351_n727# 0.29fF
C689 a_735_n727# a_351_n727# 0.05fF
C690 a_1119_n309# a_735_n309# 0.05fF
C691 a_1791_109# a_1887_109# 0.29fF
C692 a_n1857_n309# a_n1857_109# 0.01fF
C693 a_1599_109# a_1215_109# 0.05fF
C694 a_n513_n309# a_n225_n309# 0.06fF
C695 a_n129_n309# a_n321_n309# 0.11fF
C696 a_543_527# a_543_109# 0.01fF
C697 a_n993_n727# a_n993_n309# 0.01fF
C698 a_1407_n727# a_1503_n727# 0.29fF
C699 a_n225_109# a_n33_109# 0.11fF
C700 a_255_n727# a_63_n727# 0.11fF
C701 a_639_109# a_927_109# 0.06fF
C702 a_1599_n309# a_1695_n309# 0.29fF
C703 a_n1185_n309# a_n993_n309# 0.11fF
C704 a_n225_527# a_n129_527# 0.29fF
C705 a_1215_n309# a_1503_n309# 0.06fF
C706 a_735_n309# a_927_n309# 0.11fF
C707 a_1695_n727# a_1791_n727# 0.29fF
C708 a_639_n309# a_735_n309# 0.29fF
C709 a_n513_n727# a_n705_n727# 0.11fF
C710 a_n1569_n727# a_n1281_n727# 0.06fF
C711 a_351_109# a_639_109# 0.06fF
C712 a_n1185_109# a_n1185_527# 0.01fF
C713 a_n705_527# a_n705_109# 0.01fF
C714 a_1599_109# a_1407_109# 0.11fF
C715 a_543_527# a_447_527# 0.29fF
C716 a_n417_n309# a_n225_n309# 0.11fF
C717 a_1599_n727# a_1215_n727# 0.05fF
C718 a_1311_109# a_927_109# 0.05fF
C719 a_63_n309# a_63_n727# 0.01fF
C720 a_447_n309# a_447_n727# 0.01fF
C721 a_1407_n309# a_1791_n309# 0.05fF
C722 a_n1281_527# a_n993_527# 0.06fF
C723 a_n705_n727# a_n705_n309# 0.01fF
C724 a_n417_n727# a_n801_n727# 0.05fF
C725 a_n1857_527# a_n1949_527# 0.29fF
C726 a_255_n309# a_351_n309# 0.29fF
C727 a_735_n727# a_543_n727# 0.11fF
C728 a_1791_109# a_1599_109# 0.11fF
C729 a_255_n727# a_543_n727# 0.06fF
C730 a_n417_109# a_n33_109# 0.05fF
C731 a_159_n727# a_n129_n727# 0.06fF
C732 a_n1949_n727# a_n1761_n727# 0.11fF
C733 a_927_n727# a_1023_n727# 0.29fF
C734 a_n1665_n309# a_n1665_n727# 0.01fF
C735 a_n321_109# a_63_109# 0.05fF
C736 a_255_527# a_n129_527# 0.05fF
C737 a_159_n309# a_n225_n309# 0.05fF
C738 a_n1473_n727# a_n1473_n309# 0.01fF
C739 a_1887_n727# w_n2087_n937# 0.12fF
C740 a_1791_n727# w_n2087_n937# 0.08fF
C741 a_1695_n727# w_n2087_n937# 0.06fF
C742 a_1599_n727# w_n2087_n937# 0.06fF
C743 a_1503_n727# w_n2087_n937# 0.04fF
C744 a_1407_n727# w_n2087_n937# 0.04fF
C745 a_1311_n727# w_n2087_n937# 0.04fF
C746 a_1215_n727# w_n2087_n937# 0.04fF
C747 a_1119_n727# w_n2087_n937# 0.04fF
C748 a_1023_n727# w_n2087_n937# 0.04fF
C749 a_927_n727# w_n2087_n937# 0.04fF
C750 a_831_n727# w_n2087_n937# 0.04fF
C751 a_735_n727# w_n2087_n937# 0.04fF
C752 a_639_n727# w_n2087_n937# 0.04fF
C753 a_543_n727# w_n2087_n937# 0.04fF
C754 a_447_n727# w_n2087_n937# 0.04fF
C755 a_351_n727# w_n2087_n937# 0.04fF
C756 a_255_n727# w_n2087_n937# 0.04fF
C757 a_159_n727# w_n2087_n937# 0.04fF
C758 a_63_n727# w_n2087_n937# 0.04fF
C759 a_n33_n727# w_n2087_n937# 0.04fF
C760 a_n129_n727# w_n2087_n937# 0.04fF
C761 a_n225_n727# w_n2087_n937# 0.04fF
C762 a_n321_n727# w_n2087_n937# 0.04fF
C763 a_n417_n727# w_n2087_n937# 0.04fF
C764 a_n513_n727# w_n2087_n937# 0.04fF
C765 a_n609_n727# w_n2087_n937# 0.04fF
C766 a_n705_n727# w_n2087_n937# 0.04fF
C767 a_n801_n727# w_n2087_n937# 0.04fF
C768 a_n897_n727# w_n2087_n937# 0.04fF
C769 a_n993_n727# w_n2087_n937# 0.04fF
C770 a_n1089_n727# w_n2087_n937# 0.04fF
C771 a_n1185_n727# w_n2087_n937# 0.04fF
C772 a_n1281_n727# w_n2087_n937# 0.04fF
C773 a_n1377_n727# w_n2087_n937# 0.04fF
C774 a_n1473_n727# w_n2087_n937# 0.04fF
C775 a_n1569_n727# w_n2087_n937# 0.04fF
C776 a_n1665_n727# w_n2087_n937# 0.04fF
C777 a_n1761_n727# w_n2087_n937# 0.04fF
C778 a_n1857_n727# w_n2087_n937# 0.04fF
C779 a_n1949_n727# w_n2087_n937# 0.04fF
C780 a_1887_n309# w_n2087_n937# 0.11fF
C781 a_1791_n309# w_n2087_n937# 0.07fF
C782 a_1695_n309# w_n2087_n937# 0.05fF
C783 a_1599_n309# w_n2087_n937# 0.05fF
C784 a_1503_n309# w_n2087_n937# 0.03fF
C785 a_1407_n309# w_n2087_n937# 0.03fF
C786 a_1311_n309# w_n2087_n937# 0.03fF
C787 a_1215_n309# w_n2087_n937# 0.03fF
C788 a_1119_n309# w_n2087_n937# 0.03fF
C789 a_1023_n309# w_n2087_n937# 0.03fF
C790 a_927_n309# w_n2087_n937# 0.03fF
C791 a_831_n309# w_n2087_n937# 0.03fF
C792 a_735_n309# w_n2087_n937# 0.03fF
C793 a_639_n309# w_n2087_n937# 0.03fF
C794 a_543_n309# w_n2087_n937# 0.03fF
C795 a_447_n309# w_n2087_n937# 0.03fF
C796 a_351_n309# w_n2087_n937# 0.03fF
C797 a_255_n309# w_n2087_n937# 0.03fF
C798 a_159_n309# w_n2087_n937# 0.03fF
C799 a_63_n309# w_n2087_n937# 0.03fF
C800 a_n33_n309# w_n2087_n937# 0.03fF
C801 a_n129_n309# w_n2087_n937# 0.03fF
C802 a_n225_n309# w_n2087_n937# 0.03fF
C803 a_n321_n309# w_n2087_n937# 0.03fF
C804 a_n417_n309# w_n2087_n937# 0.03fF
C805 a_n513_n309# w_n2087_n937# 0.03fF
C806 a_n609_n309# w_n2087_n937# 0.03fF
C807 a_n705_n309# w_n2087_n937# 0.03fF
C808 a_n801_n309# w_n2087_n937# 0.03fF
C809 a_n897_n309# w_n2087_n937# 0.03fF
C810 a_n993_n309# w_n2087_n937# 0.03fF
C811 a_n1089_n309# w_n2087_n937# 0.03fF
C812 a_n1185_n309# w_n2087_n937# 0.03fF
C813 a_n1281_n309# w_n2087_n937# 0.03fF
C814 a_n1377_n309# w_n2087_n937# 0.03fF
C815 a_n1473_n309# w_n2087_n937# 0.03fF
C816 a_n1569_n309# w_n2087_n937# 0.03fF
C817 a_n1665_n309# w_n2087_n937# 0.03fF
C818 a_n1761_n309# w_n2087_n937# 0.03fF
C819 a_n1857_n309# w_n2087_n937# 0.03fF
C820 a_n1949_n309# w_n2087_n937# 0.03fF
C821 a_1887_109# w_n2087_n937# 0.11fF
C822 a_1791_109# w_n2087_n937# 0.07fF
C823 a_1695_109# w_n2087_n937# 0.05fF
C824 a_1599_109# w_n2087_n937# 0.05fF
C825 a_1503_109# w_n2087_n937# 0.03fF
C826 a_1407_109# w_n2087_n937# 0.03fF
C827 a_1311_109# w_n2087_n937# 0.03fF
C828 a_1215_109# w_n2087_n937# 0.03fF
C829 a_1119_109# w_n2087_n937# 0.03fF
C830 a_1023_109# w_n2087_n937# 0.03fF
C831 a_927_109# w_n2087_n937# 0.03fF
C832 a_831_109# w_n2087_n937# 0.03fF
C833 a_735_109# w_n2087_n937# 0.03fF
C834 a_639_109# w_n2087_n937# 0.03fF
C835 a_543_109# w_n2087_n937# 0.03fF
C836 a_447_109# w_n2087_n937# 0.03fF
C837 a_351_109# w_n2087_n937# 0.03fF
C838 a_255_109# w_n2087_n937# 0.03fF
C839 a_159_109# w_n2087_n937# 0.03fF
C840 a_63_109# w_n2087_n937# 0.03fF
C841 a_n33_109# w_n2087_n937# 0.03fF
C842 a_n129_109# w_n2087_n937# 0.03fF
C843 a_n225_109# w_n2087_n937# 0.03fF
C844 a_n321_109# w_n2087_n937# 0.03fF
C845 a_n417_109# w_n2087_n937# 0.03fF
C846 a_n513_109# w_n2087_n937# 0.03fF
C847 a_n609_109# w_n2087_n937# 0.03fF
C848 a_n705_109# w_n2087_n937# 0.03fF
C849 a_n801_109# w_n2087_n937# 0.03fF
C850 a_n897_109# w_n2087_n937# 0.03fF
C851 a_n993_109# w_n2087_n937# 0.03fF
C852 a_n1089_109# w_n2087_n937# 0.03fF
C853 a_n1185_109# w_n2087_n937# 0.03fF
C854 a_n1281_109# w_n2087_n937# 0.03fF
C855 a_n1377_109# w_n2087_n937# 0.03fF
C856 a_n1473_109# w_n2087_n937# 0.03fF
C857 a_n1569_109# w_n2087_n937# 0.03fF
C858 a_n1665_109# w_n2087_n937# 0.03fF
C859 a_n1761_109# w_n2087_n937# 0.03fF
C860 a_n1857_109# w_n2087_n937# 0.03fF
C861 a_n1949_109# w_n2087_n937# 0.03fF
C862 a_1887_527# w_n2087_n937# 0.12fF
C863 a_1791_527# w_n2087_n937# 0.08fF
C864 a_1695_527# w_n2087_n937# 0.06fF
C865 a_1599_527# w_n2087_n937# 0.06fF
C866 a_1503_527# w_n2087_n937# 0.04fF
C867 a_1407_527# w_n2087_n937# 0.04fF
C868 a_1311_527# w_n2087_n937# 0.04fF
C869 a_1215_527# w_n2087_n937# 0.04fF
C870 a_1119_527# w_n2087_n937# 0.04fF
C871 a_1023_527# w_n2087_n937# 0.04fF
C872 a_927_527# w_n2087_n937# 0.04fF
C873 a_831_527# w_n2087_n937# 0.04fF
C874 a_735_527# w_n2087_n937# 0.04fF
C875 a_639_527# w_n2087_n937# 0.04fF
C876 a_543_527# w_n2087_n937# 0.04fF
C877 a_447_527# w_n2087_n937# 0.04fF
C878 a_351_527# w_n2087_n937# 0.04fF
C879 a_255_527# w_n2087_n937# 0.04fF
C880 a_159_527# w_n2087_n937# 0.04fF
C881 a_63_527# w_n2087_n937# 0.04fF
C882 a_n33_527# w_n2087_n937# 0.04fF
C883 a_n129_527# w_n2087_n937# 0.04fF
C884 a_n225_527# w_n2087_n937# 0.04fF
C885 a_n321_527# w_n2087_n937# 0.04fF
C886 a_n417_527# w_n2087_n937# 0.04fF
C887 a_n513_527# w_n2087_n937# 0.04fF
C888 a_n609_527# w_n2087_n937# 0.04fF
C889 a_n705_527# w_n2087_n937# 0.04fF
C890 a_n801_527# w_n2087_n937# 0.04fF
C891 a_n897_527# w_n2087_n937# 0.04fF
C892 a_n993_527# w_n2087_n937# 0.04fF
C893 a_n1089_527# w_n2087_n937# 0.04fF
C894 a_n1185_527# w_n2087_n937# 0.04fF
C895 a_n1281_527# w_n2087_n937# 0.04fF
C896 a_n1377_527# w_n2087_n937# 0.04fF
C897 a_n1473_527# w_n2087_n937# 0.04fF
C898 a_n1569_527# w_n2087_n937# 0.04fF
C899 a_n1665_527# w_n2087_n937# 0.04fF
C900 a_n1761_527# w_n2087_n937# 0.04fF
C901 a_n1857_527# w_n2087_n937# 0.04fF
C902 a_n1949_527# w_n2087_n937# 0.04fF
C903 a_n1905_n505# w_n2087_n937# 14.96fF
.ends

.subckt source_follower_buff_nmos w_2250_n1147# out avdd1p8 avss1p8 in m1_460_n1129#
+ iref w_2049_850# w_2250_1287# w_2250_355#
Xsky130_fd_pr__nfet_01v8_lvt_CFLRKA_0 avdd1p8 out out out out out avdd1p8 out out
+ out avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 out avdd1p8
+ avdd1p8 out avdd1p8 out out avdd1p8 out avdd1p8 out out out avdd1p8 out avdd1p8
+ out avss1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 out avdd1p8 out avdd1p8
+ avdd1p8 avdd1p8 out out out out avdd1p8 out out out avdd1p8 out avdd1p8 avdd1p8
+ avdd1p8 avdd1p8 out out out avdd1p8 avdd1p8 out out out out avdd1p8 out out avdd1p8
+ avdd1p8 in avdd1p8 avdd1p8 avdd1p8 out out avdd1p8 out sky130_fd_pr__nfet_01v8_lvt_CFLRKA
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_0 m1_460_n1129# iref iref iref m1_460_n1129# m1_460_n1129#
+ avss1p8 m1_460_n1129# iref sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_1 avss1p8 m1_460_n1129# m1_460_n1129# iref avss1p8
+ avss1p8 avss1p8 avss1p8 m1_460_n1129# sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_CAF2P9_0 out out avss1p8 out avss1p8 out out out out
+ avss1p8 out out avss1p8 out out out avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 out
+ avss1p8 out out avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 iref out avss1p8
+ out out out avss1p8 avss1p8 avss1p8 out out avss1p8 avss1p8 out avss1p8 avss1p8
+ out out avss1p8 out out out out out out out avss1p8 avss1p8 avss1p8 out out out
+ out out out avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 out avss1p8 avss1p8
+ avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 out out avss1p8 avss1p8 avss1p8
+ avss1p8 avss1p8 avss1p8 avss1p8 out out out out out out avss1p8 avss1p8 out avss1p8
+ out out out out out avss1p8 out out out avss1p8 avss1p8 out avss1p8 avss1p8 avss1p8
+ avss1p8 out avss1p8 out avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 out out
+ out avss1p8 avss1p8 out avss1p8 avss1p8 avss1p8 out out out out avss1p8 out avss1p8
+ avss1p8 out out out out out avss1p8 avss1p8 out avss1p8 out avss1p8 out out avss1p8
+ avss1p8 avss1p8 avss1p8 avss1p8 out out out avss1p8 avss1p8 out sky130_fd_pr__nfet_01v8_lvt_CAF2P9
C0 iref m1_460_n1129# 2.64fF
C1 out in 10.03fF
C2 iref in 0.11fF
C3 out iref 22.08fF
C4 avdd1p8 in 2.17fF
C5 avdd1p8 out 9.98fF
C6 iref avss1p8 18.70fF
C7 in avss1p8 -31.17fF
C8 out avss1p8 -28.37fF
C9 m1_460_n1129# avss1p8 2.61fF
C10 avdd1p8 avss1p8 2.63fF
.ends

.subckt source_follower_buff_diff outn VSUBS avdd1p8 inp source_follower_buff_pmos_0/m1_957_828#
+ iref1 outp iref2 iref3 iref4 source_follower_buff_nmos_1/m1_460_n1129# source_follower_buff_pmos_1/m1_957_828#
+ source_follower_buff_nmos_0/in source_follower_buff_nmos_0/m1_460_n1129# source_follower_buff_nmos_1/in
+ source_follower_buff_nmos_0/w_2250_355# inn
Xsource_follower_buff_pmos_0 source_follower_buff_pmos_0/m1_957_828# inn VSUBS avdd1p8
+ source_follower_buff_nmos_0/in iref3 source_follower_buff_pmos
Xsource_follower_buff_pmos_1 source_follower_buff_pmos_1/m1_957_828# inp VSUBS avdd1p8
+ source_follower_buff_nmos_1/in iref1 source_follower_buff_pmos
Xsource_follower_buff_nmos_0 source_follower_buff_nmos_0/w_2250_n1147# outn avdd1p8
+ VSUBS source_follower_buff_nmos_0/in source_follower_buff_nmos_0/m1_460_n1129# iref4
+ source_follower_buff_nmos_0/w_2049_850# source_follower_buff_nmos_0/w_2250_1287#
+ source_follower_buff_nmos_0/w_2250_355# source_follower_buff_nmos
Xsource_follower_buff_nmos_1 source_follower_buff_nmos_1/w_2250_n1147# outp avdd1p8
+ VSUBS source_follower_buff_nmos_1/in source_follower_buff_nmos_1/m1_460_n1129# iref2
+ source_follower_buff_nmos_1/w_2049_850# source_follower_buff_nmos_1/w_2250_1287#
+ source_follower_buff_nmos_1/w_2250_355# source_follower_buff_nmos
C0 source_follower_buff_nmos_1/in avdd1p8 0.63fF
C1 inp avdd1p8 0.07fF
C2 outn avdd1p8 0.18fF
C3 outp source_follower_buff_nmos_1/w_2250_n1147# 0.09fF
C4 inp source_follower_buff_pmos_1/m1_957_828# 0.08fF
C5 inn source_follower_buff_nmos_0/in -0.25fF
C6 source_follower_buff_nmos_0/w_2049_850# avdd1p8 0.16fF
C7 outn source_follower_buff_nmos_0/in 0.11fF
C8 inp source_follower_buff_nmos_1/in -0.25fF
C9 inn source_follower_buff_pmos_0/m1_957_828# 0.08fF
C10 outp source_follower_buff_nmos_1/in 0.11fF
C11 source_follower_buff_nmos_0/w_2250_1287# avdd1p8 0.18fF
C12 iref3 inn 0.01fF
C13 inn avdd1p8 0.07fF
C14 source_follower_buff_nmos_0/in avdd1p8 0.63fF
C15 inp iref1 0.01fF
C16 iref2 VSUBS 11.84fF
C17 source_follower_buff_nmos_1/in VSUBS -32.98fF
C18 outp VSUBS 0.56fF
C19 source_follower_buff_nmos_1/m1_460_n1129# VSUBS 1.47fF
C20 iref4 VSUBS 12.04fF
C21 source_follower_buff_nmos_0/in VSUBS -32.98fF
C22 outn VSUBS 2.12fF
C23 source_follower_buff_nmos_0/m1_460_n1129# VSUBS 1.50fF
C24 avdd1p8 VSUBS 35.96fF
C25 inp VSUBS 2.70fF
C26 source_follower_buff_pmos_1/m1_957_828# VSUBS -35.44fF
C27 iref1 VSUBS 3.02fF
C28 inn VSUBS 4.09fF
C29 source_follower_buff_pmos_0/m1_957_828# VSUBS -35.44fF
C30 iref3 VSUBS 3.13fF
.ends

.subckt res_amp_top avss1p8 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_3/in
+ avdd1p8 iref0 res_amp_lin_prog_0/res_amp_lin_0/a_3747_261# iref1 res_amp_lin_prog_0/res_amp_lin_0/vp
+ res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/out iref2 res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/in1
+ res_amp_lin_prog_0/outn iref3 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1384_n363#
+ res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/out source_follower_buff_diff_0/source_follower_buff_pmos_0/m1_957_828#
+ delay_reg0 iref4 res_amp_lin_prog_0/outp res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/in
+ res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/inverter_min_1/in res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinB
+ inn source_follower_buff_diff_0/source_follower_buff_pmos_1/m1_957_828# inp res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_511_801#
+ res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/sel_b res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_12/inverter_min_1/in
+ res_amp_lin_prog_0/res_amp_lin_0/clk res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinA
+ res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/DinA delay_reg2 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_5/out
+ res_amp_lin_prog_0/outp_cap iref_reg0 res_amp_lin_prog_0/clk res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinB
+ source_follower_buff_diff_0/source_follower_buff_nmos_1/in res_amp_lin_prog_0/res_amp_lin_0/vctrl
+ res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_2/inverter_min_1/in res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinA
+ res_amp_sync_v2_0/clkp iref_reg1 source_follower_buff_diff_0/source_follower_buff_nmos_0/in
+ res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/out iref_reg2 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_964_n363#
+ res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_10/inverter_min_1/in res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/out
+ res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/sel_b res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/out
+ res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/m1_21_n341# res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_7/inverter_min_1/in
+ delay_reg1 outn source_follower_buff_diff_0/source_follower_buff_nmos_1/m1_460_n1129#
+ outp clkn res_amp_sync_v2_0/rst
Xres_amp_sync_v2_0 avdd1p8 res_amp_sync_v2_0/DFlipFlop_4/Q avss1p8 clkn res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/m1_657_280#
+ res_amp_sync_v2_0/DFlipFlop_4/nQ res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/nD res_amp_sync_v2_0/DFlipFlop_3/latch_diff_0/D
+ res_amp_sync_v2_0/DFlipFlop_3/Q res_amp_sync_v2_0/DFlipFlop_3/D res_amp_sync_v2_0/DFlipFlop_4/D
+ res_amp_sync_v2_0/DFlipFlop_1/D res_amp_sync_v2_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/D res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/nD
+ res_amp_sync_v2_0/DFlipFlop_4/clock_inverter_0/inverter_cp_x1_2/in res_amp_sync_v2_0/DFlipFlop_4/latch_diff_0/D
+ res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/D res_amp_lin_prog_0/clk res_amp_sync_v2_0/DFlipFlop_3/nQ
+ res_amp_sync_v2_0/clkp res_amp_sync_v2_0/rst res_amp_sync_v2
Xres_amp_lin_prog_0 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/out res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_964_n363#
+ delay_reg2 avdd1p8 inp res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinA
+ res_amp_lin_prog_0/res_amp_lin_0/vctrl res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/out
+ res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_511_801# res_amp_lin_prog_0/res_amp_lin_0/clk
+ res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/in1 res_amp_lin_prog_0/outp_cap
+ avss1p8 res_amp_lin_prog_0/outn_cap res_amp_lin_prog_0/clk res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/sel_b
+ delay_reg0 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinA res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinB
+ res_amp_lin_prog_0/outn res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/DinA
+ res_amp_lin_prog_0/outp res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_5/out
+ res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_2/inverter_min_1/in res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinB
+ iref_reg0 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/inverter_min_1/in
+ iref_reg1 iref_reg2 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1384_n363# res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_3/in
+ res_amp_lin_prog_0/res_amp_lin_0/vp res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/m1_21_n341#
+ res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/out res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/out
+ res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_12/inverter_min_1/in iref0
+ res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_7/inverter_min_1/in res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_n356_n363#
+ res_amp_lin_prog_0/res_amp_lin_0/a_3747_261# delay_reg1 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/in
+ inn res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/out res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1996_n363#
+ res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_10/inverter_min_1/in res_amp_lin_prog_0/inverter_min_x4_0/out
+ res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/sel_b res_amp_sync_v2_0/rst
+ res_amp_lin_prog
Xsky130_fd_pr__cap_mim_m3_1_U5ZKVF_0 avss1p8 avss1p8 res_amp_lin_prog_0/outp_cap sky130_fd_pr__cap_mim_m3_1_U5ZKVF
Xsky130_fd_pr__cap_mim_m3_1_U5ZKVF_1 avss1p8 avss1p8 res_amp_lin_prog_0/outn_cap sky130_fd_pr__cap_mim_m3_1_U5ZKVF
Xsource_follower_buff_diff_0 outn avss1p8 avdd1p8 res_amp_lin_prog_0/outp_cap source_follower_buff_diff_0/source_follower_buff_pmos_0/m1_957_828#
+ iref1 outp iref2 iref3 iref4 source_follower_buff_diff_0/source_follower_buff_nmos_1/m1_460_n1129#
+ source_follower_buff_diff_0/source_follower_buff_pmos_1/m1_957_828# source_follower_buff_diff_0/source_follower_buff_nmos_0/in
+ source_follower_buff_diff_0/source_follower_buff_nmos_0/m1_460_n1129# source_follower_buff_diff_0/source_follower_buff_nmos_1/in
+ source_follower_buff_diff_0/source_follower_buff_nmos_0/w_2250_355# res_amp_lin_prog_0/outn_cap
+ source_follower_buff_diff
C0 res_amp_sync_v2_0/DFlipFlop_3/D res_amp_lin_prog_0/clk 0.07fF
C1 avdd1p8 source_follower_buff_diff_0/source_follower_buff_pmos_1/m1_957_828# 0.02fF
C2 res_amp_lin_prog_0/clk res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/nD 0.25fF
C3 res_amp_lin_prog_0/res_amp_lin_0/vctrl iref0 -0.03fF
C4 delay_reg1 avdd1p8 0.04fF
C5 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1996_n363# avdd1p8 1.10fF
C6 res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/D res_amp_lin_prog_0/clk 0.23fF
C7 avdd1p8 res_amp_lin_prog_0/clk 9.77fF
C8 avdd1p8 clkn 0.74fF
C9 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/out delay_reg2 0.03fF
C10 inp res_amp_sync_v2_0/rst 0.09fF
C11 avdd1p8 delay_reg2 0.08fF
C12 res_amp_sync_v2_0/DFlipFlop_4/Q res_amp_lin_prog_0/clk 0.44fF
C13 avdd1p8 source_follower_buff_diff_0/source_follower_buff_nmos_1/in 0.40fF
C14 res_amp_sync_v2_0/clkp clkn 0.06fF
C15 res_amp_lin_prog_0/clk res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/nD 0.28fF
C16 res_amp_sync_v2_0/rst avdd1p8 0.80fF
C17 delay_reg0 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/out 0.04fF
C18 res_amp_sync_v2_0/rst res_amp_lin_prog_0/outp_cap 0.13fF
C19 avdd1p8 res_amp_sync_v2_0/DFlipFlop_3/D 0.89fF
C20 iref3 source_follower_buff_diff_0/source_follower_buff_pmos_0/m1_957_828# 0.10fF
C21 inp avdd1p8 0.46fF
C22 avdd1p8 res_amp_sync_v2_0/DFlipFlop_1/D 0.29fF
C23 res_amp_lin_prog_0/clk res_amp_sync_v2_0/DFlipFlop_3/Q 0.25fF
C24 res_amp_lin_prog_0/clk res_amp_sync_v2_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in 0.48fF
C25 res_amp_sync_v2_0/DFlipFlop_3/nQ res_amp_lin_prog_0/clk 0.20fF
C26 res_amp_sync_v2_0/rst res_amp_lin_prog_0/outn_cap 0.06fF
C27 outn source_follower_buff_diff_0/source_follower_buff_nmos_0/w_2250_355# 0.15fF
C28 avdd1p8 outp 0.31fF
C29 iref_reg1 avdd1p8 0.05fF
C30 res_amp_sync_v2_0/clkp avdd1p8 1.19fF
C31 res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/m1_657_280# res_amp_lin_prog_0/clk 0.06fF
C32 source_follower_buff_diff_0/source_follower_buff_pmos_0/m1_957_828# avdd1p8 0.02fF
C33 avdd1p8 source_follower_buff_diff_0/source_follower_buff_nmos_0/in 0.39fF
C34 res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/D res_amp_lin_prog_0/clk 0.20fF
C35 res_amp_sync_v2_0/DFlipFlop_4/latch_diff_0/D res_amp_lin_prog_0/clk 0.47fF
C36 iref0 avdd1p8 -0.63fF
C37 iref2 source_follower_buff_diff_0/source_follower_buff_nmos_1/m1_460_n1129# 0.12fF
C38 outn avdd1p8 0.30fF
C39 iref0 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1384_n363# 0.02fF
C40 iref4 source_follower_buff_diff_0/source_follower_buff_nmos_0/m1_460_n1129# 0.13fF
C41 res_amp_sync_v2_0/DFlipFlop_3/latch_diff_0/D res_amp_lin_prog_0/clk 0.47fF
C42 iref1 source_follower_buff_diff_0/source_follower_buff_pmos_1/m1_957_828# 0.10fF
C43 res_amp_sync_v2_0/DFlipFlop_4/D res_amp_lin_prog_0/clk 0.08fF
C44 res_amp_sync_v2_0/rst inn 0.09fF
C45 res_amp_sync_v2_0/DFlipFlop_4/nQ res_amp_lin_prog_0/clk 0.22fF
C46 res_amp_lin_prog_0/clk clkn 0.07fF
C47 inp inn 1.68fF
C48 delay_reg1 delay_reg2 0.23fF
C49 res_amp_lin_prog_0/res_amp_lin_0/vctrl avdd1p8 0.03fF
C50 avdd1p8 iref_reg2 -0.57fF
C51 avdd1p8 inn 0.46fF
C52 res_amp_sync_v2_0/DFlipFlop_4/clock_inverter_0/inverter_cp_x1_2/in res_amp_lin_prog_0/clk 0.48fF
C53 iref2 avss1p8 12.17fF
C54 source_follower_buff_diff_0/source_follower_buff_nmos_1/in avss1p8 -32.88fF
C55 outp avss1p8 -1.74fF
C56 source_follower_buff_diff_0/source_follower_buff_nmos_1/m1_460_n1129# avss1p8 1.82fF
C57 iref4 avss1p8 12.36fF
C58 source_follower_buff_diff_0/source_follower_buff_nmos_0/in avss1p8 -32.87fF
C59 source_follower_buff_diff_0/source_follower_buff_nmos_0/w_2250_355# avss1p8 0.08fF
C60 outn avss1p8 -1.13fF
C61 source_follower_buff_diff_0/source_follower_buff_nmos_0/m1_460_n1129# avss1p8 1.84fF
C62 source_follower_buff_diff_0/source_follower_buff_pmos_1/m1_957_828# avss1p8 -35.44fF
C63 iref1 avss1p8 3.33fF
C64 source_follower_buff_diff_0/source_follower_buff_pmos_0/m1_957_828# avss1p8 -35.44fF
C65 iref3 avss1p8 3.02fF
C66 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_511_801# avss1p8 -1.87fF
C67 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1384_n363# avss1p8 0.47fF
C68 iref_reg1 avss1p8 0.41fF
C69 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_448_n363# avss1p8 -1.10fF
C70 res_amp_lin_prog_0/res_amp_lin_0/vctrl avss1p8 -1.99fF
C71 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1996_n363# avss1p8 -2.18fF
C72 iref_reg2 avss1p8 0.06fF
C73 iref_reg0 avss1p8 -0.21fF
C74 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_964_n363# avss1p8 -1.03fF
C75 res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_n356_n363# avss1p8 0.55fF
C76 iref0 avss1p8 0.37fF
C77 res_amp_lin_prog_0/outn avss1p8 1.55fF
C78 inp avss1p8 0.21fF
C79 res_amp_lin_prog_0/outp avss1p8 -4.89fF
C80 res_amp_lin_prog_0/res_amp_lin_0/vp avss1p8 -4.89fF
C81 inn avss1p8 -6.68fF
C82 res_amp_lin_prog_0/res_amp_lin_0/a_3747_261# avss1p8 -0.95fF
C83 res_amp_lin_prog_0/outn_cap avss1p8 1.00fF
C84 res_amp_lin_prog_0/inverter_min_x4_0/out avss1p8 4.87fF
C85 res_amp_lin_prog_0/res_amp_lin_0/clk avss1p8 4.30fF
C86 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_7/in avss1p8 1.07fF
C87 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinA avss1p8 -0.04fF
C88 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_7/inverter_min_1/in avss1p8 1.03fF
C89 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_6/inverter_min_1/in avss1p8 1.03fF
C90 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_5/in avss1p8 1.07fF
C91 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_5/inverter_min_1/in avss1p8 1.03fF
C92 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_4/inverter_min_1/in avss1p8 1.03fF
C93 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_3/in avss1p8 1.07fF
C94 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_3/inverter_min_1/in avss1p8 1.03fF
C95 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_1/in avss1p8 1.07fF
C96 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_1/inverter_min_1/in avss1p8 1.03fF
C97 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_2/inverter_min_1/in avss1p8 1.03fF
C98 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_0/inverter_min_1/in avss1p8 1.04fF
C99 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/in avss1p8 1.07fF
C100 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinB avss1p8 -7.88fF
C101 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/inverter_min_1/in avss1p8 1.03fF
C102 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_12/inverter_min_1/in avss1p8 1.03fF
C103 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_11/in avss1p8 1.07fF
C104 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_11/inverter_min_1/in avss1p8 1.03fF
C105 res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/m1_21_n341# avss1p8 0.72fF
C106 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_10/inverter_min_1/in avss1p8 1.03fF
C107 res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/in1 avss1p8 1.54fF
C108 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_6/sel_b avss1p8 2.03fF
C109 delay_reg0 avss1p8 2.90fF
C110 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_5/out avss1p8 -1.67fF
C111 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_5/sel_b avss1p8 2.03fF
C112 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinA avss1p8 -2.58fF
C113 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/out avss1p8 -2.25fF
C114 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/sel_b avss1p8 2.03fF
C115 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/out avss1p8 -2.69fF
C116 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinB avss1p8 -4.96fF
C117 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/sel_b avss1p8 2.03fF
C118 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/out avss1p8 -4.71fF
C119 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/sel_b avss1p8 2.03fF
C120 delay_reg1 avss1p8 3.97fF
C121 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/DinA avss1p8 0.63fF
C122 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/out avss1p8 -2.49fF
C123 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/DinB avss1p8 -3.92fF
C124 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/sel_b avss1p8 2.03fF
C125 delay_reg2 avss1p8 11.33fF
C126 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/out avss1p8 -0.27fF
C127 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/DinB avss1p8 -0.97fF
C128 res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/sel_b avss1p8 2.04fF
C129 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_9/in avss1p8 1.07fF
C130 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_9/inverter_min_1/in avss1p8 1.03fF
C131 res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_8/inverter_min_1/in avss1p8 1.03fF
C132 res_amp_lin_prog_0/outp_cap avss1p8 -6.67fF
C133 res_amp_sync_v2_0/nand_logic_1/m1_21_n341# avss1p8 0.72fF
C134 res_amp_sync_v2_0/nand_logic_0/m1_21_n341# avss1p8 0.72fF
C135 res_amp_lin_prog_0/clk avss1p8 -6.90fF
C136 res_amp_sync_v2_0/inverter_min_x4_4/out avss1p8 5.85fF
C137 res_amp_sync_v2_0/rst avss1p8 -3.03fF
C138 res_amp_sync_v2_0/nand_logic_1/out avss1p8 1.70fF
C139 res_amp_sync_v2_0/DFlipFlop_4/Q avss1p8 -2.08fF
C140 res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/m1_657_280# avss1p8 0.57fF
C141 res_amp_sync_v2_0/DFlipFlop_4/nQ avss1p8 0.48fF
C142 res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/D avss1p8 -1.73fF
C143 res_amp_sync_v2_0/DFlipFlop_4/latch_diff_0/m1_657_280# avss1p8 0.57fF
C144 res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/nD avss1p8 0.57fF
C145 res_amp_sync_v2_0/DFlipFlop_4/clock_inverter_0/inverter_cp_x1_2/in avss1p8 1.86fF
C146 res_amp_sync_v2_0/DFlipFlop_4/latch_diff_0/D avss1p8 0.96fF
C147 res_amp_sync_v2_0/DFlipFlop_4/clock_inverter_0/inverter_cp_x1_0/out avss1p8 1.76fF
C148 res_amp_sync_v2_0/DFlipFlop_4/D avss1p8 1.83fF
C149 res_amp_sync_v2_0/DFlipFlop_4/latch_diff_0/nD avss1p8 1.14fF
C150 res_amp_sync_v2_0/nand_logic_0/out avss1p8 1.20fF
C151 res_amp_sync_v2_0/DFlipFlop_3/Q avss1p8 -2.94fF
C152 res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/m1_657_280# avss1p8 0.57fF
C153 clkn avss1p8 -7.50fF
C154 res_amp_sync_v2_0/DFlipFlop_3/nQ avss1p8 0.48fF
C155 res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/D avss1p8 -1.73fF
C156 res_amp_sync_v2_0/DFlipFlop_3/latch_diff_0/m1_657_280# avss1p8 0.57fF
C157 res_amp_sync_v2_0/clkp avss1p8 -28.00fF
C158 res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/nD avss1p8 0.57fF
C159 res_amp_sync_v2_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in avss1p8 1.86fF
C160 res_amp_sync_v2_0/DFlipFlop_3/latch_diff_0/D avss1p8 0.96fF
C161 res_amp_sync_v2_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out avss1p8 1.76fF
C162 res_amp_sync_v2_0/DFlipFlop_3/D avss1p8 1.33fF
C163 avdd1p8 avss1p8 415.30fF
C164 res_amp_sync_v2_0/DFlipFlop_3/latch_diff_0/nD avss1p8 1.14fF
C165 res_amp_sync_v2_0/DFlipFlop_2/Q avss1p8 -1.08fF
C166 res_amp_sync_v2_0/DFlipFlop_2/latch_diff_1/m1_657_280# avss1p8 0.57fF
C167 res_amp_sync_v2_0/DFlipFlop_2/nQ avss1p8 0.48fF
C168 res_amp_sync_v2_0/DFlipFlop_2/latch_diff_1/D avss1p8 -1.73fF
C169 res_amp_sync_v2_0/DFlipFlop_2/latch_diff_0/m1_657_280# avss1p8 0.57fF
C170 res_amp_sync_v2_0/DFlipFlop_2/latch_diff_1/nD avss1p8 0.57fF
C171 res_amp_sync_v2_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in avss1p8 1.86fF
C172 res_amp_sync_v2_0/DFlipFlop_2/latch_diff_0/D avss1p8 0.96fF
C173 res_amp_sync_v2_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out avss1p8 1.76fF
C174 res_amp_sync_v2_0/DFlipFlop_2/D avss1p8 -0.38fF
C175 res_amp_sync_v2_0/DFlipFlop_2/latch_diff_0/nD avss1p8 1.14fF
C176 res_amp_sync_v2_0/DFlipFlop_1/latch_diff_1/m1_657_280# avss1p8 0.57fF
C177 res_amp_sync_v2_0/DFlipFlop_1/nQ avss1p8 0.48fF
C178 res_amp_sync_v2_0/DFlipFlop_1/latch_diff_1/D avss1p8 -1.73fF
C179 res_amp_sync_v2_0/DFlipFlop_1/latch_diff_0/m1_657_280# avss1p8 0.57fF
C180 res_amp_sync_v2_0/DFlipFlop_1/latch_diff_1/nD avss1p8 0.57fF
C181 res_amp_sync_v2_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in avss1p8 1.86fF
C182 res_amp_sync_v2_0/DFlipFlop_1/latch_diff_0/D avss1p8 0.96fF
C183 res_amp_sync_v2_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out avss1p8 1.76fF
C184 res_amp_sync_v2_0/DFlipFlop_1/D avss1p8 -1.02fF
C185 res_amp_sync_v2_0/DFlipFlop_1/latch_diff_0/nD avss1p8 1.14fF
C186 res_amp_sync_v2_0/DFlipFlop_0/Q avss1p8 -4.73fF
C187 res_amp_sync_v2_0/DFlipFlop_0/latch_diff_1/m1_657_280# avss1p8 0.57fF
C188 res_amp_sync_v2_0/DFlipFlop_0/nQ avss1p8 0.48fF
C189 res_amp_sync_v2_0/DFlipFlop_0/latch_diff_1/D avss1p8 -1.73fF
C190 res_amp_sync_v2_0/DFlipFlop_0/latch_diff_0/m1_657_280# avss1p8 0.57fF
C191 res_amp_sync_v2_0/DFlipFlop_0/latch_diff_1/nD avss1p8 0.57fF
C192 res_amp_sync_v2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in avss1p8 1.86fF
C193 res_amp_sync_v2_0/DFlipFlop_0/latch_diff_0/D avss1p8 0.96fF
C194 res_amp_sync_v2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out avss1p8 1.76fF
C195 res_amp_sync_v2_0/DFlipFlop_0/latch_diff_0/nD avss1p8 1.14fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4ML9WA VSUBS a_429_n486# w_n2457_n634# a_887_n486#
+ a_n29_n486# a_1345_n486# a_n2261_n512# a_1803_n486# a_n487_n486# a_n945_n486# a_n2319_n486#
+ a_n1403_n486# a_2261_n486# a_n1861_n486#
X0 a_2261_n486# a_n2261_n512# a_1803_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X1 a_n945_n486# a_n2261_n512# a_n1403_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X2 a_429_n486# a_n2261_n512# a_n29_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X3 a_1803_n486# a_n2261_n512# a_1345_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X4 a_887_n486# a_n2261_n512# a_429_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X5 a_n487_n486# a_n2261_n512# a_n945_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X6 a_n1403_n486# a_n2261_n512# a_n1861_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X7 a_n1861_n486# a_n2261_n512# a_n2319_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X8 a_n29_n486# a_n2261_n512# a_n487_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X9 a_1345_n486# a_n2261_n512# a_887_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
C0 w_n2457_n634# a_n1861_n486# 0.02fF
C1 a_n945_n486# w_n2457_n634# 0.02fF
C2 w_n2457_n634# a_n487_n486# 0.02fF
C3 w_n2457_n634# a_n1403_n486# 0.02fF
C4 a_429_n486# w_n2457_n634# 0.02fF
C5 a_n29_n486# w_n2457_n634# 0.02fF
C6 w_n2457_n634# a_2261_n486# 0.02fF
C7 a_n2319_n486# w_n2457_n634# 0.02fF
C8 w_n2457_n634# a_887_n486# 0.02fF
C9 w_n2457_n634# a_1345_n486# 0.02fF
C10 a_1803_n486# w_n2457_n634# 0.02fF
C11 a_2261_n486# VSUBS 0.03fF
C12 a_1803_n486# VSUBS 0.03fF
C13 a_1345_n486# VSUBS 0.03fF
C14 a_887_n486# VSUBS 0.03fF
C15 a_429_n486# VSUBS 0.03fF
C16 a_n29_n486# VSUBS 0.03fF
C17 a_n487_n486# VSUBS 0.03fF
C18 a_n945_n486# VSUBS 0.03fF
C19 a_n1403_n486# VSUBS 0.03fF
C20 a_n1861_n486# VSUBS 0.03fF
C21 a_n2319_n486# VSUBS 0.03fF
C22 a_n2261_n512# VSUBS 4.27fF
C23 w_n2457_n634# VSUBS 21.34fF
.ends

.subckt sky130_fd_pr__nfet_01v8_YCGG98 a_n1041_n75# a_n561_n75# a_1167_n75# a_303_n75#
+ a_687_n75# a_n849_n75# a_n369_n75# a_975_n75# a_111_n75# a_495_n75# a_n1137_n75#
+ a_n657_n75# a_n177_n75# a_783_n75# a_n945_n75# a_n465_n75# a_207_n75# a_1071_n75#
+ a_591_n75# a_15_n75# a_n753_n75# w_n1367_n285# a_n273_n75# a_879_n75# a_399_n75#
+ a_n1229_n75# a_n81_n75# a_n1167_n101#
X0 a_207_n75# a_n1167_n101# a_111_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_303_n75# a_n1167_n101# a_207_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_399_n75# a_n1167_n101# a_303_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_495_n75# a_n1167_n101# a_399_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_591_n75# a_n1167_n101# a_495_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_783_n75# a_n1167_n101# a_687_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_687_n75# a_n1167_n101# a_591_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_879_n75# a_n1167_n101# a_783_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_975_n75# a_n1167_n101# a_879_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_n1041_n75# a_n1167_n101# a_n1137_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_n1137_n75# a_n1167_n101# a_n1229_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n561_n75# a_n1167_n101# a_n657_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_1071_n75# a_n1167_n101# a_975_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n945_n75# a_n1167_n101# a_n1041_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n753_n75# a_n1167_n101# a_n849_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n657_n75# a_n1167_n101# a_n753_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n465_n75# a_n1167_n101# a_n561_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n369_n75# a_n1167_n101# a_n465_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_1167_n75# a_n1167_n101# a_1071_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n849_n75# a_n1167_n101# a_n945_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X20 a_15_n75# a_n1167_n101# a_n81_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X21 a_n81_n75# a_n1167_n101# a_n177_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X22 a_111_n75# a_n1167_n101# a_15_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X23 a_n273_n75# a_n1167_n101# a_n369_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X24 a_n177_n75# a_n1167_n101# a_n273_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
C0 a_n561_n75# a_n369_n75# 0.08fF
C1 a_495_n75# a_687_n75# 0.08fF
C2 a_n753_n75# a_n369_n75# 0.03fF
C3 a_399_n75# a_495_n75# 0.22fF
C4 a_n1041_n75# a_n1137_n75# 0.22fF
C5 a_n849_n75# a_n1229_n75# 0.03fF
C6 a_n273_n75# a_n657_n75# 0.03fF
C7 a_n465_n75# a_n657_n75# 0.08fF
C8 a_n753_n75# a_n1137_n75# 0.03fF
C9 a_399_n75# a_111_n75# 0.05fF
C10 a_n1041_n75# a_n753_n75# 0.05fF
C11 a_n753_n75# a_n561_n75# 0.08fF
C12 a_n849_n75# a_n1137_n75# 0.05fF
C13 a_15_n75# a_n273_n75# 0.05fF
C14 a_111_n75# a_495_n75# 0.03fF
C15 a_15_n75# a_n81_n75# 0.22fF
C16 a_n1041_n75# a_n849_n75# 0.08fF
C17 a_15_n75# a_n177_n75# 0.08fF
C18 a_n561_n75# a_n849_n75# 0.05fF
C19 a_n753_n75# a_n849_n75# 0.22fF
C20 a_n273_n75# a_n369_n75# 0.22fF
C21 a_n81_n75# a_n369_n75# 0.05fF
C22 a_591_n75# a_207_n75# 0.03fF
C23 a_n465_n75# a_n369_n75# 0.22fF
C24 a_n177_n75# a_n369_n75# 0.08fF
C25 a_15_n75# a_207_n75# 0.08fF
C26 a_975_n75# a_783_n75# 0.08fF
C27 a_n561_n75# a_n273_n75# 0.05fF
C28 a_n657_n75# a_n945_n75# 0.05fF
C29 a_591_n75# a_303_n75# 0.05fF
C30 a_n465_n75# a_n561_n75# 0.22fF
C31 a_n561_n75# a_n177_n75# 0.03fF
C32 a_15_n75# a_303_n75# 0.05fF
C33 a_975_n75# a_1167_n75# 0.08fF
C34 a_n465_n75# a_n753_n75# 0.05fF
C35 a_1167_n75# a_783_n75# 0.03fF
C36 a_111_n75# a_n273_n75# 0.03fF
C37 a_399_n75# a_207_n75# 0.08fF
C38 a_111_n75# a_n81_n75# 0.08fF
C39 a_111_n75# a_n177_n75# 0.05fF
C40 a_n465_n75# a_n849_n75# 0.03fF
C41 a_975_n75# a_1071_n75# 0.22fF
C42 a_207_n75# a_495_n75# 0.05fF
C43 a_975_n75# a_591_n75# 0.03fF
C44 a_1071_n75# a_783_n75# 0.05fF
C45 a_303_n75# a_687_n75# 0.03fF
C46 a_591_n75# a_783_n75# 0.08fF
C47 a_975_n75# a_879_n75# 0.22fF
C48 a_n945_n75# a_n1229_n75# 0.05fF
C49 a_399_n75# a_303_n75# 0.22fF
C50 a_879_n75# a_783_n75# 0.22fF
C51 a_111_n75# a_207_n75# 0.22fF
C52 a_1071_n75# a_1167_n75# 0.22fF
C53 a_495_n75# a_303_n75# 0.08fF
C54 a_1167_n75# a_879_n75# 0.05fF
C55 a_n1137_n75# a_n945_n75# 0.08fF
C56 a_n81_n75# a_n273_n75# 0.08fF
C57 a_n465_n75# a_n273_n75# 0.08fF
C58 a_975_n75# a_687_n75# 0.05fF
C59 a_n177_n75# a_n273_n75# 0.22fF
C60 a_n1041_n75# a_n945_n75# 0.22fF
C61 a_n465_n75# a_n81_n75# 0.03fF
C62 a_n561_n75# a_n945_n75# 0.03fF
C63 a_783_n75# a_687_n75# 0.22fF
C64 a_n81_n75# a_n177_n75# 0.22fF
C65 a_n465_n75# a_n177_n75# 0.05fF
C66 a_111_n75# a_303_n75# 0.08fF
C67 a_399_n75# a_783_n75# 0.03fF
C68 a_1071_n75# a_879_n75# 0.08fF
C69 a_n753_n75# a_n945_n75# 0.08fF
C70 a_591_n75# a_879_n75# 0.05fF
C71 a_n657_n75# a_n369_n75# 0.05fF
C72 a_783_n75# a_495_n75# 0.05fF
C73 a_n849_n75# a_n945_n75# 0.22fF
C74 a_207_n75# a_n81_n75# 0.05fF
C75 a_207_n75# a_n177_n75# 0.03fF
C76 a_1071_n75# a_687_n75# 0.03fF
C77 a_15_n75# a_n369_n75# 0.03fF
C78 a_591_n75# a_687_n75# 0.22fF
C79 a_n1041_n75# a_n657_n75# 0.03fF
C80 a_n561_n75# a_n657_n75# 0.22fF
C81 a_879_n75# a_687_n75# 0.08fF
C82 a_399_n75# a_591_n75# 0.08fF
C83 a_399_n75# a_15_n75# 0.03fF
C84 a_n81_n75# a_303_n75# 0.03fF
C85 a_n753_n75# a_n657_n75# 0.22fF
C86 a_591_n75# a_495_n75# 0.22fF
C87 a_879_n75# a_495_n75# 0.03fF
C88 a_n849_n75# a_n657_n75# 0.08fF
C89 a_n1137_n75# a_n1229_n75# 0.22fF
C90 a_399_n75# a_687_n75# 0.05fF
C91 a_207_n75# a_303_n75# 0.22fF
C92 a_n1041_n75# a_n1229_n75# 0.08fF
C93 a_15_n75# a_111_n75# 0.22fF
C94 a_1167_n75# w_n1367_n285# 0.10fF
C95 a_1071_n75# w_n1367_n285# 0.07fF
C96 a_975_n75# w_n1367_n285# 0.06fF
C97 a_879_n75# w_n1367_n285# 0.05fF
C98 a_783_n75# w_n1367_n285# 0.04fF
C99 a_687_n75# w_n1367_n285# 0.04fF
C100 a_591_n75# w_n1367_n285# 0.04fF
C101 a_495_n75# w_n1367_n285# 0.04fF
C102 a_399_n75# w_n1367_n285# 0.04fF
C103 a_303_n75# w_n1367_n285# 0.04fF
C104 a_207_n75# w_n1367_n285# 0.04fF
C105 a_111_n75# w_n1367_n285# 0.04fF
C106 a_15_n75# w_n1367_n285# 0.04fF
C107 a_n81_n75# w_n1367_n285# 0.04fF
C108 a_n177_n75# w_n1367_n285# 0.04fF
C109 a_n273_n75# w_n1367_n285# 0.04fF
C110 a_n369_n75# w_n1367_n285# 0.04fF
C111 a_n465_n75# w_n1367_n285# 0.04fF
C112 a_n561_n75# w_n1367_n285# 0.04fF
C113 a_n657_n75# w_n1367_n285# 0.04fF
C114 a_n753_n75# w_n1367_n285# 0.04fF
C115 a_n849_n75# w_n1367_n285# 0.04fF
C116 a_n945_n75# w_n1367_n285# 0.04fF
C117 a_n1041_n75# w_n1367_n285# 0.04fF
C118 a_n1137_n75# w_n1367_n285# 0.04fF
C119 a_n1229_n75# w_n1367_n285# 0.04fF
C120 a_n1167_n101# w_n1367_n285# 2.55fF
.ends

.subckt sky130_fd_pr__nfet_01v8_MUHGM9 a_33_n101# a_n129_n75# a_735_n75# a_255_n75#
+ a_n417_n75# a_n989_n75# a_63_n75# a_543_n75# a_n705_n75# a_n225_n75# a_n33_n75#
+ a_831_n75# a_351_n75# a_n927_n101# a_n513_n75# a_n897_n75# w_n1127_n285# a_639_n75#
+ a_159_n75# a_n801_n75# a_n321_n75# a_927_n75# a_447_n75# a_n609_n75#
X0 a_63_n75# a_33_n101# a_n33_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_927_n75# a_33_n101# a_831_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_n33_n75# a_n927_n101# a_n129_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_159_n75# a_33_n101# a_63_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_255_n75# a_33_n101# a_159_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_351_n75# a_33_n101# a_255_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_447_n75# a_33_n101# a_351_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_543_n75# a_33_n101# a_447_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_735_n75# a_33_n101# a_639_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_831_n75# a_33_n101# a_735_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_639_n75# a_33_n101# a_543_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n321_n75# a_n927_n101# a_n417_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_n801_n75# a_n927_n101# a_n897_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n705_n75# a_n927_n101# a_n801_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n513_n75# a_n927_n101# a_n609_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n417_n75# a_n927_n101# a_n513_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n225_n75# a_n927_n101# a_n321_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n129_n75# a_n927_n101# a_n225_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_n897_n75# a_n927_n101# a_n989_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n609_n75# a_n927_n101# a_n705_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
C0 a_n225_n75# a_n513_n75# 0.05fF
C1 a_n225_n75# a_63_n75# 0.05fF
C2 a_255_n75# a_639_n75# 0.03fF
C3 a_447_n75# a_735_n75# 0.05fF
C4 a_n225_n75# a_159_n75# 0.03fF
C5 a_447_n75# a_639_n75# 0.08fF
C6 a_n321_n75# a_n609_n75# 0.05fF
C7 a_255_n75# a_543_n75# 0.05fF
C8 a_n801_n75# a_n609_n75# 0.08fF
C9 a_n321_n75# a_n129_n75# 0.08fF
C10 a_n321_n75# a_n705_n75# 0.03fF
C11 a_447_n75# a_543_n75# 0.22fF
C12 a_n801_n75# a_n705_n75# 0.22fF
C13 a_n321_n75# a_n417_n75# 0.22fF
C14 a_543_n75# a_159_n75# 0.03fF
C15 a_n33_n75# a_351_n75# 0.03fF
C16 a_n801_n75# a_n417_n75# 0.03fF
C17 a_927_n75# a_831_n75# 0.22fF
C18 a_n609_n75# a_n705_n75# 0.22fF
C19 a_n33_n75# a_n321_n75# 0.05fF
C20 a_n417_n75# a_n609_n75# 0.08fF
C21 a_n417_n75# a_n129_n75# 0.05fF
C22 a_735_n75# a_639_n75# 0.22fF
C23 a_n417_n75# a_n705_n75# 0.05fF
C24 a_n801_n75# a_n989_n75# 0.08fF
C25 a_n33_n75# a_n129_n75# 0.22fF
C26 a_n989_n75# a_n609_n75# 0.03fF
C27 a_543_n75# a_735_n75# 0.08fF
C28 a_543_n75# a_639_n75# 0.22fF
C29 a_n33_n75# a_n417_n75# 0.03fF
C30 a_n989_n75# a_n705_n75# 0.05fF
C31 a_255_n75# a_351_n75# 0.22fF
C32 a_351_n75# a_63_n75# 0.05fF
C33 a_n801_n75# a_n897_n75# 0.22fF
C34 a_n321_n75# a_n513_n75# 0.08fF
C35 a_447_n75# a_351_n75# 0.22fF
C36 a_n801_n75# a_n513_n75# 0.05fF
C37 a_n927_n101# a_33_n101# 0.08fF
C38 a_n321_n75# a_63_n75# 0.03fF
C39 a_351_n75# a_159_n75# 0.08fF
C40 a_447_n75# a_831_n75# 0.03fF
C41 a_n609_n75# a_n897_n75# 0.05fF
C42 a_n513_n75# a_n609_n75# 0.22fF
C43 a_n897_n75# a_n705_n75# 0.08fF
C44 a_n513_n75# a_n129_n75# 0.03fF
C45 a_n513_n75# a_n705_n75# 0.08fF
C46 a_255_n75# a_n129_n75# 0.03fF
C47 a_63_n75# a_n129_n75# 0.08fF
C48 a_n513_n75# a_n417_n75# 0.22fF
C49 a_n129_n75# a_159_n75# 0.05fF
C50 a_735_n75# a_351_n75# 0.03fF
C51 a_351_n75# a_639_n75# 0.05fF
C52 a_n989_n75# a_n897_n75# 0.22fF
C53 a_255_n75# a_n33_n75# 0.05fF
C54 a_n33_n75# a_63_n75# 0.22fF
C55 a_n225_n75# a_n321_n75# 0.22fF
C56 a_735_n75# a_831_n75# 0.22fF
C57 a_831_n75# a_639_n75# 0.08fF
C58 a_n33_n75# a_159_n75# 0.08fF
C59 a_543_n75# a_351_n75# 0.08fF
C60 a_n225_n75# a_n609_n75# 0.03fF
C61 a_n225_n75# a_n129_n75# 0.22fF
C62 a_543_n75# a_831_n75# 0.05fF
C63 a_n225_n75# a_n417_n75# 0.08fF
C64 a_927_n75# a_735_n75# 0.08fF
C65 a_n513_n75# a_n897_n75# 0.03fF
C66 a_927_n75# a_639_n75# 0.05fF
C67 a_n225_n75# a_n33_n75# 0.08fF
C68 a_255_n75# a_63_n75# 0.08fF
C69 a_927_n75# a_543_n75# 0.03fF
C70 a_447_n75# a_255_n75# 0.08fF
C71 a_447_n75# a_63_n75# 0.03fF
C72 a_255_n75# a_159_n75# 0.22fF
C73 a_63_n75# a_159_n75# 0.22fF
C74 a_447_n75# a_159_n75# 0.05fF
C75 a_927_n75# w_n1127_n285# 0.04fF
C76 a_831_n75# w_n1127_n285# 0.04fF
C77 a_735_n75# w_n1127_n285# 0.04fF
C78 a_639_n75# w_n1127_n285# 0.04fF
C79 a_543_n75# w_n1127_n285# 0.04fF
C80 a_447_n75# w_n1127_n285# 0.04fF
C81 a_351_n75# w_n1127_n285# 0.04fF
C82 a_255_n75# w_n1127_n285# 0.04fF
C83 a_159_n75# w_n1127_n285# 0.04fF
C84 a_63_n75# w_n1127_n285# 0.04fF
C85 a_n33_n75# w_n1127_n285# 0.04fF
C86 a_n129_n75# w_n1127_n285# 0.04fF
C87 a_n225_n75# w_n1127_n285# 0.04fF
C88 a_n321_n75# w_n1127_n285# 0.04fF
C89 a_n417_n75# w_n1127_n285# 0.04fF
C90 a_n513_n75# w_n1127_n285# 0.04fF
C91 a_n609_n75# w_n1127_n285# 0.04fF
C92 a_n705_n75# w_n1127_n285# 0.04fF
C93 a_n801_n75# w_n1127_n285# 0.04fF
C94 a_n897_n75# w_n1127_n285# 0.04fF
C95 a_n989_n75# w_n1127_n285# 0.04fF
C96 a_33_n101# w_n1127_n285# 0.99fF
C97 a_n927_n101# w_n1127_n285# 0.99fF
.ends

.subckt sky130_fd_pr__pfet_01v8_NKZXKB VSUBS a_33_n247# a_n801_n150# a_n417_n150#
+ a_351_n150# a_255_n150# a_n705_n150# a_n609_n150# a_159_n150# a_543_n150# a_447_n150#
+ a_831_n150# a_n897_n150# a_n33_n150# a_735_n150# a_n927_n247# a_639_n150# a_n321_n150#
+ a_927_n150# a_n225_n150# a_63_n150# a_n989_n150# a_n513_n150# a_n129_n150# w_n1127_n369#
X0 a_n513_n150# a_n927_n247# a_n609_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_63_n150# a_33_n247# a_n33_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_735_n150# a_33_n247# a_639_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n801_n150# a_n927_n247# a_n897_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n927_n247# a_n225_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n927_n247# a_n513_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_639_n150# a_33_n247# a_543_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n705_n150# a_n927_n247# a_n801_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n33_n150# a_n927_n247# a_n129_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_351_n150# a_33_n247# a_255_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_n609_n150# a_n927_n247# a_n705_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n897_n150# a_n927_n247# a_n989_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_927_n150# a_33_n247# a_831_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_255_n150# a_33_n247# a_159_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n321_n150# a_n927_n247# a_n417_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_543_n150# a_33_n247# a_447_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_831_n150# a_33_n247# a_735_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_159_n150# a_33_n247# a_63_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_n225_n150# a_n927_n247# a_n321_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_447_n150# a_33_n247# a_351_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n417_n150# a_n705_n150# 0.10fF
C1 a_n609_n150# a_n513_n150# 0.43fF
C2 a_63_n150# a_n225_n150# 0.10fF
C3 a_n609_n150# a_n225_n150# 0.07fF
C4 a_735_n150# a_927_n150# 0.16fF
C5 a_n897_n150# a_n513_n150# 0.07fF
C6 a_351_n150# a_735_n150# 0.07fF
C7 a_n609_n150# a_n989_n150# 0.07fF
C8 a_n927_n247# a_33_n247# 0.09fF
C9 a_n417_n150# a_n513_n150# 0.43fF
C10 a_159_n150# a_543_n150# 0.07fF
C11 a_351_n150# a_n33_n150# 0.07fF
C12 a_735_n150# a_447_n150# 0.10fF
C13 a_n417_n150# a_n225_n150# 0.16fF
C14 a_n897_n150# a_n989_n150# 0.43fF
C15 a_255_n150# a_543_n150# 0.10fF
C16 a_639_n150# a_831_n150# 0.16fF
C17 a_639_n150# a_543_n150# 0.43fF
C18 a_n897_n150# a_n609_n150# 0.10fF
C19 a_n33_n150# a_n225_n150# 0.16fF
C20 a_n417_n150# a_n609_n150# 0.16fF
C21 a_63_n150# a_n33_n150# 0.43fF
C22 a_n705_n150# a_n321_n150# 0.07fF
C23 a_n705_n150# a_n801_n150# 0.43fF
C24 a_159_n150# a_351_n150# 0.16fF
C25 a_255_n150# a_351_n150# 0.43fF
C26 a_159_n150# a_447_n150# 0.10fF
C27 a_n129_n150# a_n513_n150# 0.07fF
C28 a_639_n150# a_927_n150# 0.10fF
C29 a_n417_n150# a_n33_n150# 0.07fF
C30 a_n129_n150# a_n225_n150# 0.43fF
C31 a_639_n150# a_351_n150# 0.10fF
C32 a_543_n150# a_831_n150# 0.10fF
C33 a_255_n150# a_447_n150# 0.16fF
C34 a_n513_n150# a_n321_n150# 0.16fF
C35 a_n513_n150# a_n801_n150# 0.10fF
C36 a_159_n150# a_n225_n150# 0.07fF
C37 a_n225_n150# a_n321_n150# 0.43fF
C38 a_639_n150# a_447_n150# 0.16fF
C39 a_n129_n150# a_63_n150# 0.16fF
C40 a_n989_n150# a_n801_n150# 0.16fF
C41 a_159_n150# a_63_n150# 0.43fF
C42 a_63_n150# a_n321_n150# 0.07fF
C43 a_n609_n150# a_n321_n150# 0.10fF
C44 a_n609_n150# a_n801_n150# 0.16fF
C45 a_255_n150# a_63_n150# 0.16fF
C46 a_n417_n150# a_n129_n150# 0.10fF
C47 a_n897_n150# a_n801_n150# 0.43fF
C48 a_n417_n150# a_n321_n150# 0.43fF
C49 a_n417_n150# a_n801_n150# 0.07fF
C50 a_927_n150# a_831_n150# 0.43fF
C51 a_543_n150# a_927_n150# 0.07fF
C52 a_351_n150# a_543_n150# 0.16fF
C53 a_n129_n150# a_n33_n150# 0.43fF
C54 a_447_n150# a_831_n150# 0.07fF
C55 a_543_n150# a_447_n150# 0.43fF
C56 a_159_n150# a_n33_n150# 0.16fF
C57 a_n33_n150# a_n321_n150# 0.10fF
C58 a_639_n150# a_735_n150# 0.43fF
C59 a_255_n150# a_n33_n150# 0.10fF
C60 a_n705_n150# a_n513_n150# 0.16fF
C61 a_159_n150# a_n129_n150# 0.10fF
C62 a_n129_n150# a_n321_n150# 0.16fF
C63 a_351_n150# a_447_n150# 0.43fF
C64 a_255_n150# a_n129_n150# 0.07fF
C65 a_735_n150# a_831_n150# 0.43fF
C66 a_543_n150# a_735_n150# 0.16fF
C67 a_255_n150# a_159_n150# 0.43fF
C68 a_n989_n150# a_n705_n150# 0.10fF
C69 a_n609_n150# a_n705_n150# 0.43fF
C70 a_639_n150# a_255_n150# 0.07fF
C71 a_n225_n150# a_n513_n150# 0.10fF
C72 a_351_n150# a_63_n150# 0.10fF
C73 a_n897_n150# a_n705_n150# 0.16fF
C74 a_63_n150# a_447_n150# 0.07fF
C75 a_927_n150# VSUBS 0.03fF
C76 a_831_n150# VSUBS 0.03fF
C77 a_735_n150# VSUBS 0.03fF
C78 a_639_n150# VSUBS 0.03fF
C79 a_543_n150# VSUBS 0.03fF
C80 a_447_n150# VSUBS 0.03fF
C81 a_351_n150# VSUBS 0.03fF
C82 a_255_n150# VSUBS 0.03fF
C83 a_159_n150# VSUBS 0.03fF
C84 a_63_n150# VSUBS 0.03fF
C85 a_n33_n150# VSUBS 0.03fF
C86 a_n129_n150# VSUBS 0.03fF
C87 a_n225_n150# VSUBS 0.03fF
C88 a_n321_n150# VSUBS 0.03fF
C89 a_n417_n150# VSUBS 0.03fF
C90 a_n513_n150# VSUBS 0.03fF
C91 a_n609_n150# VSUBS 0.03fF
C92 a_n705_n150# VSUBS 0.03fF
C93 a_n801_n150# VSUBS 0.03fF
C94 a_n897_n150# VSUBS 0.03fF
C95 a_n989_n150# VSUBS 0.03fF
C96 a_33_n247# VSUBS 1.04fF
C97 a_n927_n247# VSUBS 1.04fF
C98 w_n1127_n369# VSUBS 6.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_8GRULZ a_n1761_n132# a_1045_n44# a_n1461_n44# a_n1103_n44#
+ a_n29_n44# a_n387_n44# a_1761_n44# a_n1819_n44# a_1403_n44# a_687_n44# w_n1957_n254#
+ a_329_n44# a_n745_n44#
X0 a_329_n44# a_n1761_n132# a_n29_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X1 a_1761_n44# a_n1761_n132# a_1403_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X2 a_n745_n44# a_n1761_n132# a_n1103_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X3 a_1045_n44# a_n1761_n132# a_687_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X4 a_n29_n44# a_n1761_n132# a_n387_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X5 a_n1103_n44# a_n1761_n132# a_n1461_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X6 a_n387_n44# a_n1761_n132# a_n745_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X7 a_687_n44# a_n1761_n132# a_329_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X8 a_1403_n44# a_n1761_n132# a_1045_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X9 a_n1461_n44# a_n1761_n132# a_n1819_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
C0 a_1761_n44# a_1403_n44# 0.04fF
C1 a_329_n44# a_n29_n44# 0.04fF
C2 a_n29_n44# a_n387_n44# 0.04fF
C3 a_329_n44# a_687_n44# 0.04fF
C4 a_n745_n44# a_n1103_n44# 0.04fF
C5 a_n1819_n44# a_n1461_n44# 0.04fF
C6 a_1045_n44# a_1403_n44# 0.04fF
C7 a_687_n44# a_1045_n44# 0.04fF
C8 a_n745_n44# a_n387_n44# 0.04fF
C9 a_n1461_n44# a_n1103_n44# 0.04fF
C10 a_1761_n44# w_n1957_n254# 0.04fF
C11 a_1403_n44# w_n1957_n254# 0.04fF
C12 a_1045_n44# w_n1957_n254# 0.04fF
C13 a_687_n44# w_n1957_n254# 0.04fF
C14 a_329_n44# w_n1957_n254# 0.04fF
C15 a_n29_n44# w_n1957_n254# 0.04fF
C16 a_n387_n44# w_n1957_n254# 0.04fF
C17 a_n745_n44# w_n1957_n254# 0.04fF
C18 a_n1103_n44# w_n1957_n254# 0.04fF
C19 a_n1461_n44# w_n1957_n254# 0.04fF
C20 a_n1819_n44# w_n1957_n254# 0.04fF
C21 a_n1761_n132# w_n1957_n254# 3.23fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ND88ZC VSUBS a_303_n150# a_n753_n150# a_n369_n150#
+ w_n1367_n369# a_207_n150# a_n657_n150# a_591_n150# a_n1229_n150# a_n945_n150# a_495_n150#
+ a_n1041_n150# a_n849_n150# a_n81_n150# a_399_n150# a_783_n150# a_1071_n150# a_687_n150#
+ a_975_n150# a_n1137_n150# a_n273_n150# a_111_n150# a_879_n150# a_n177_n150# a_n561_n150#
+ a_15_n150# a_1167_n150# a_n1167_n247# a_n465_n150#
X0 a_n1137_n150# a_n1167_n247# a_n1229_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_495_n150# a_n1167_n247# a_399_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n561_n150# a_n1167_n247# a_n657_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_111_n150# a_n1167_n247# a_15_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_783_n150# a_n1167_n247# a_687_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_1071_n150# a_n1167_n247# a_975_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_399_n150# a_n1167_n247# a_303_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n465_n150# a_n1167_n247# a_n561_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_687_n150# a_n1167_n247# a_591_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n753_n150# a_n1167_n247# a_n849_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_975_n150# a_n1167_n247# a_879_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n81_n150# a_n1167_n247# a_n177_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_15_n150# a_n1167_n247# a_n81_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_n1041_n150# a_n1167_n247# a_n1137_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n369_n150# a_n1167_n247# a_n465_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_n657_n150# a_n1167_n247# a_n753_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_879_n150# a_n1167_n247# a_783_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_n945_n150# a_n1167_n247# a_n1041_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_1167_n150# a_n1167_n247# a_1071_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_303_n150# a_n1167_n247# a_207_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X20 a_n273_n150# a_n1167_n247# a_n369_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X21 a_591_n150# a_n1167_n247# a_495_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X22 a_n849_n150# a_n1167_n247# a_n945_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_207_n150# a_n1167_n247# a_111_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X24 a_n177_n150# a_n1167_n247# a_n273_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n945_n150# a_n561_n150# 0.07fF
C1 a_303_n150# a_15_n150# 0.10fF
C2 a_n753_n150# a_n945_n150# 0.16fF
C3 a_n1137_n150# a_n1229_n150# 0.43fF
C4 a_n465_n150# a_n273_n150# 0.16fF
C5 a_1167_n150# a_879_n150# 0.10fF
C6 a_n177_n150# a_n369_n150# 0.16fF
C7 a_783_n150# a_1167_n150# 0.07fF
C8 w_n1367_n369# a_1071_n150# 0.07fF
C9 a_n465_n150# a_n81_n150# 0.07fF
C10 a_495_n150# a_207_n150# 0.10fF
C11 a_783_n150# a_399_n150# 0.07fF
C12 a_207_n150# a_591_n150# 0.07fF
C13 a_399_n150# a_687_n150# 0.10fF
C14 a_n657_n150# a_n561_n150# 0.43fF
C15 a_n849_n150# a_n1137_n150# 0.10fF
C16 a_495_n150# a_399_n150# 0.43fF
C17 a_n657_n150# a_n753_n150# 0.43fF
C18 a_399_n150# a_591_n150# 0.16fF
C19 a_n177_n150# a_n273_n150# 0.43fF
C20 a_n1041_n150# a_n1229_n150# 0.16fF
C21 a_n177_n150# a_207_n150# 0.07fF
C22 a_n753_n150# a_n561_n150# 0.16fF
C23 a_303_n150# a_687_n150# 0.07fF
C24 a_n657_n150# a_n465_n150# 0.16fF
C25 a_n945_n150# a_n1229_n150# 0.10fF
C26 a_111_n150# a_n273_n150# 0.07fF
C27 a_975_n150# a_879_n150# 0.43fF
C28 a_303_n150# a_495_n150# 0.16fF
C29 a_111_n150# a_207_n150# 0.43fF
C30 a_303_n150# a_591_n150# 0.10fF
C31 a_n177_n150# a_n81_n150# 0.43fF
C32 a_n465_n150# a_n561_n150# 0.43fF
C33 a_n465_n150# a_n753_n150# 0.10fF
C34 a_111_n150# a_399_n150# 0.10fF
C35 a_783_n150# a_975_n150# 0.16fF
C36 a_975_n150# a_687_n150# 0.10fF
C37 a_n849_n150# a_n1041_n150# 0.16fF
C38 a_111_n150# a_n81_n150# 0.16fF
C39 a_1071_n150# a_1167_n150# 0.43fF
C40 a_n177_n150# a_15_n150# 0.16fF
C41 a_975_n150# a_591_n150# 0.07fF
C42 w_n1367_n369# a_1167_n150# 0.14fF
C43 a_n849_n150# a_n945_n150# 0.43fF
C44 a_783_n150# a_879_n150# 0.43fF
C45 a_303_n150# a_111_n150# 0.16fF
C46 a_879_n150# a_687_n150# 0.16fF
C47 a_111_n150# a_15_n150# 0.43fF
C48 a_n1041_n150# a_n1137_n150# 0.43fF
C49 a_495_n150# a_879_n150# 0.07fF
C50 a_879_n150# a_591_n150# 0.10fF
C51 a_n177_n150# a_n561_n150# 0.07fF
C52 a_n945_n150# a_n1137_n150# 0.16fF
C53 a_783_n150# a_687_n150# 0.43fF
C54 a_n369_n150# a_n273_n150# 0.43fF
C55 a_783_n150# a_495_n150# 0.10fF
C56 a_495_n150# a_687_n150# 0.16fF
C57 a_783_n150# a_591_n150# 0.16fF
C58 a_591_n150# a_687_n150# 0.43fF
C59 a_n465_n150# a_n177_n150# 0.10fF
C60 a_n849_n150# a_n657_n150# 0.16fF
C61 a_495_n150# a_591_n150# 0.43fF
C62 a_n81_n150# a_n369_n150# 0.10fF
C63 a_n849_n150# a_n561_n150# 0.10fF
C64 a_1071_n150# a_975_n150# 0.43fF
C65 a_n849_n150# a_n753_n150# 0.43fF
C66 w_n1367_n369# a_975_n150# 0.05fF
C67 a_399_n150# a_207_n150# 0.16fF
C68 a_n1041_n150# a_n945_n150# 0.43fF
C69 a_1071_n150# a_879_n150# 0.16fF
C70 a_15_n150# a_n369_n150# 0.07fF
C71 a_n849_n150# a_n465_n150# 0.07fF
C72 a_n81_n150# a_n273_n150# 0.16fF
C73 a_495_n150# a_111_n150# 0.07fF
C74 w_n1367_n369# a_879_n150# 0.04fF
C75 a_n753_n150# a_n1137_n150# 0.07fF
C76 a_n81_n150# a_207_n150# 0.10fF
C77 a_n657_n150# a_n369_n150# 0.10fF
C78 a_783_n150# a_1071_n150# 0.10fF
C79 a_303_n150# a_207_n150# 0.43fF
C80 a_n561_n150# a_n369_n150# 0.16fF
C81 a_1071_n150# a_687_n150# 0.07fF
C82 a_n753_n150# a_n369_n150# 0.07fF
C83 a_15_n150# a_n273_n150# 0.10fF
C84 a_n177_n150# a_111_n150# 0.10fF
C85 a_15_n150# a_207_n150# 0.16fF
C86 a_303_n150# a_399_n150# 0.43fF
C87 a_n657_n150# a_n273_n150# 0.07fF
C88 a_n657_n150# a_n1041_n150# 0.07fF
C89 a_15_n150# a_399_n150# 0.07fF
C90 a_303_n150# a_n81_n150# 0.07fF
C91 a_n465_n150# a_n369_n150# 0.43fF
C92 a_n849_n150# a_n1229_n150# 0.07fF
C93 a_n561_n150# a_n273_n150# 0.10fF
C94 a_n81_n150# a_15_n150# 0.43fF
C95 a_975_n150# a_1167_n150# 0.16fF
C96 a_n657_n150# a_n945_n150# 0.10fF
C97 a_n1041_n150# a_n753_n150# 0.10fF
C98 a_1167_n150# VSUBS 0.03fF
C99 a_1071_n150# VSUBS 0.03fF
C100 a_975_n150# VSUBS 0.03fF
C101 a_879_n150# VSUBS 0.03fF
C102 a_783_n150# VSUBS 0.03fF
C103 a_687_n150# VSUBS 0.03fF
C104 a_591_n150# VSUBS 0.03fF
C105 a_495_n150# VSUBS 0.03fF
C106 a_399_n150# VSUBS 0.03fF
C107 a_303_n150# VSUBS 0.03fF
C108 a_207_n150# VSUBS 0.03fF
C109 a_111_n150# VSUBS 0.03fF
C110 a_15_n150# VSUBS 0.03fF
C111 a_n81_n150# VSUBS 0.03fF
C112 a_n177_n150# VSUBS 0.03fF
C113 a_n273_n150# VSUBS 0.03fF
C114 a_n369_n150# VSUBS 0.03fF
C115 a_n465_n150# VSUBS 0.03fF
C116 a_n561_n150# VSUBS 0.03fF
C117 a_n657_n150# VSUBS 0.03fF
C118 a_n753_n150# VSUBS 0.03fF
C119 a_n849_n150# VSUBS 0.03fF
C120 a_n945_n150# VSUBS 0.03fF
C121 a_n1041_n150# VSUBS 0.03fF
C122 a_n1137_n150# VSUBS 0.03fF
C123 a_n1229_n150# VSUBS 0.03fF
C124 a_n1167_n247# VSUBS 2.63fF
C125 w_n1367_n369# VSUBS 7.85fF
.ends

.subckt charge_pump vss pswitch nswitch out vdd biasp nUp Down w_2544_775# iref nDown
+ Up w_1008_774# w_6648_570#
Xsky130_fd_pr__pfet_01v8_4ML9WA_0 vss pswitch vdd pswitch pswitch pswitch nUp pswitch
+ pswitch pswitch pswitch pswitch pswitch pswitch sky130_fd_pr__pfet_01v8_4ML9WA
Xsky130_fd_pr__nfet_01v8_YCGG98_0 vss out out vss vss vss out out vss vss out vss
+ out out out vss out vss out out out vss vss vss out vss vss nswitch sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_1 iref vss vss iref iref iref vss vss iref iref vss
+ iref vss vss vss iref vss iref vss vss vss vss iref iref vss iref iref iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_2 biasp vss vss biasp biasp biasp vss vss biasp biasp
+ vss biasp vss vss vss biasp vss biasp vss vss vss vss biasp biasp vss biasp biasp
+ iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_MUHGM9_0 nDown iref nswitch vss nswitch nswitch vss nswitch
+ iref nswitch nswitch vss nswitch Down iref iref vss vss nswitch nswitch iref nswitch
+ vss nswitch sky130_fd_pr__nfet_01v8_MUHGM9
Xsky130_fd_pr__pfet_01v8_NKZXKB_0 vss Up pswitch pswitch pswitch vdd biasp pswitch
+ pswitch pswitch vdd vdd biasp pswitch pswitch nUp vdd biasp pswitch pswitch vdd
+ pswitch biasp biasp vdd sky130_fd_pr__pfet_01v8_NKZXKB
Xsky130_fd_pr__nfet_01v8_8GRULZ_0 Down nswitch nswitch nswitch nswitch nswitch nswitch
+ nswitch nswitch nswitch vss nswitch nswitch sky130_fd_pr__nfet_01v8_8GRULZ
Xsky130_fd_pr__pfet_01v8_ND88ZC_0 vss vdd out out vdd out vdd out vdd out vdd vdd
+ vdd vdd out out vdd vdd out out vdd vdd vdd out out out out pswitch vdd sky130_fd_pr__pfet_01v8_ND88ZC
Xsky130_fd_pr__pfet_01v8_ND88ZC_1 vss biasp vdd vdd vdd vdd biasp vdd biasp vdd biasp
+ biasp biasp biasp vdd vdd biasp biasp vdd vdd biasp biasp biasp vdd vdd vdd vdd
+ biasp biasp sky130_fd_pr__pfet_01v8_ND88ZC
C0 nUp Up 0.15fF
C1 nswitch pswitch 0.06fF
C2 out pswitch 4.91fF
C3 vdd biasp 2.64fF
C4 nswitch biasp 0.03fF
C5 nswitch iref 1.91fF
C6 Down nDown 0.13fF
C7 nUp Down 0.25fF
C8 pswitch biasp 3.11fF
C9 pswitch Up 0.70fF
C10 nswitch nDown 0.31fF
C11 out nUp 0.31fF
C12 pswitch nUp 5.66fF
C13 nswitch vdd 0.07fF
C14 vdd out 6.66fF
C15 iref biasp 0.80fF
C16 vdd pswitch 3.98fF
C17 nswitch Down 2.27fF
C18 nswitch out 1.28fF
C19 vdd vss 35.71fF
C20 Down vss 4.77fF
C21 Up vss 1.17fF
C22 nswitch vss 6.39fF
C23 nDown vss 1.11fF
C24 biasp vss 8.73fF
C25 iref vss 10.12fF
C26 out vss -3.49fF
C27 pswitch vss 3.45fF
C28 nUp vss 5.85fF
.ends

.subckt sky130_fd_pr__nfet_01v8_5RJ8EK a_n33_n42# a_33_n68# w_n263_n252# a_n63_n68#
+ a_n125_n42# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n125_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_63_n42# a_n125_n42# 0.05fF
C1 a_n125_n42# a_n33_n42# 0.12fF
C2 a_n63_n68# a_33_n68# 0.02fF
C3 a_63_n42# a_n33_n42# 0.12fF
C4 a_63_n42# w_n263_n252# 0.09fF
C5 a_n33_n42# w_n263_n252# 0.07fF
C6 a_n125_n42# w_n263_n252# 0.09fF
C7 a_33_n68# w_n263_n252# 0.05fF
C8 a_n63_n68# w_n263_n252# 0.05fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ZPB9BB VSUBS a_n63_n110# a_33_n110# a_n125_n84# a_63_n84#
+ w_n263_n303# a_n33_n84#
X0 a_63_n84# a_33_n110# a_n33_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_n33_n84# a_n63_n110# a_n125_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_63_n84# a_n33_n84# 0.24fF
C1 a_63_n84# a_n125_n84# 0.09fF
C2 a_63_n84# w_n263_n303# 0.10fF
C3 a_n33_n84# a_n125_n84# 0.24fF
C4 a_n33_n84# w_n263_n303# 0.07fF
C5 a_33_n110# a_n63_n110# 0.02fF
C6 w_n263_n303# a_n125_n84# 0.10fF
C7 a_63_n84# VSUBS 0.03fF
C8 a_n33_n84# VSUBS 0.03fF
C9 a_n125_n84# VSUBS 0.03fF
C10 a_33_n110# VSUBS 0.05fF
C11 a_n63_n110# VSUBS 0.05fF
C12 w_n263_n303# VSUBS 1.74fF
.ends

.subckt inverter_min_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_5RJ8EK_0 vss in vss in out out sky130_fd_pr__nfet_01v8_5RJ8EK
Xsky130_fd_pr__pfet_01v8_ZPB9BB_0 vss in in out out vdd vdd sky130_fd_pr__pfet_01v8_ZPB9BB
C0 out vdd 0.15fF
C1 out in 0.30fF
C2 in vdd 0.01fF
C3 vdd vss 2.93fF
C4 out vss 0.66fF
C5 in vss 0.72fF
.ends

.subckt div_by_2 vss vdd nout_div clock_inverter_0/inverter_cp_x1_2/in CLK_2 nCLK_2
+ o1 CLK out_div o2 clock_inverter_0/inverter_cp_x1_0/out
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vss vdd DFlipFlop_0/latch_diff_1/D
+ DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in nout_div DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_0/nD
+ out_div DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/latch_diff_1/m1_657_280# nout_div
+ DFlipFlop_0/latch_diff_0/D DFlipFlop_0/CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
Xinverter_min_x4_1 vdd o2 vss nCLK_2 inverter_min_x4
Xinverter_min_x4_0 vdd o1 vss CLK_2 inverter_min_x4
Xclock_inverter_0 vss clock_inverter_0/inverter_cp_x1_2/in CLK vdd clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_0/CLK DFlipFlop_0/nCLK clock_inverter
Xinverter_min_x2_0 nout_div o2 vss vdd inverter_min_x2
Xinverter_min_x2_1 out_div o1 vss vdd inverter_min_x2
C0 DFlipFlop_0/latch_diff_1/m1_657_280# nout_div 0.21fF
C1 out_div vdd 0.03fF
C2 DFlipFlop_0/latch_diff_1/D nout_div 0.64fF
C3 DFlipFlop_0/latch_diff_0/nD nout_div 0.07fF
C4 vdd DFlipFlop_0/CLK 0.40fF
C5 DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/CLK 0.11fF
C6 DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_0/D 0.13fF
C7 DFlipFlop_0/latch_diff_0/m1_657_280# nout_div 0.24fF
C8 o1 out_div 0.01fF
C9 DFlipFlop_0/latch_diff_1/D DFlipFlop_0/CLK -0.48fF
C10 DFlipFlop_0/CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.29fF
C11 o2 vdd 0.14fF
C12 DFlipFlop_0/latch_diff_0/nD DFlipFlop_0/CLK 0.12fF
C13 out_div nout_div 0.22fF
C14 DFlipFlop_0/nCLK vdd 0.30fF
C15 DFlipFlop_0/CLK nout_div 0.42fF
C16 o2 DFlipFlop_0/latch_diff_1/m1_657_280# 0.02fF
C17 vdd CLK_2 0.08fF
C18 clock_inverter_0/inverter_cp_x1_0/out vdd 0.10fF
C19 DFlipFlop_0/latch_diff_0/m1_657_280# DFlipFlop_0/CLK 0.26fF
C20 DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/nCLK -0.09fF
C21 DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_1/m1_657_280# 0.26fF
C22 o2 nCLK_2 0.11fF
C23 DFlipFlop_0/latch_diff_0/D nout_div 0.09fF
C24 vdd DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.03fF
C25 DFlipFlop_0/nCLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.46fF
C26 DFlipFlop_0/latch_diff_1/D DFlipFlop_0/nCLK 0.08fF
C27 vdd DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C28 vdd nCLK_2 0.08fF
C29 o1 vdd 0.14fF
C30 vdd nout_div 0.16fF
C31 DFlipFlop_0/nCLK nout_div 0.43fF
C32 o1 CLK_2 0.11fF
C33 o1 DFlipFlop_0/latch_diff_1/m1_657_280# 0.02fF
C34 DFlipFlop_0/latch_diff_1/nD nout_div 1.18fF
C35 clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C36 DFlipFlop_0/CLK vss 1.03fF
C37 clock_inverter_0/inverter_cp_x1_0/out vss 1.85fF
C38 CLK vss 3.27fF
C39 DFlipFlop_0/nCLK vss 1.76fF
C40 CLK_2 vss 1.08fF
C41 o1 vss 2.21fF
C42 nCLK_2 vss 1.08fF
C43 o2 vss 2.21fF
C44 out_div vss -0.77fF
C45 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.63fF
C46 DFlipFlop_0/latch_diff_1/D vss -1.72fF
C47 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C48 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C49 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.89fF
C50 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C51 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.80fF
C52 nout_div vss 4.41fF
C53 vdd vss 64.43fF
C54 DFlipFlop_0/latch_diff_0/nD vss 1.14fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MACBVW VSUBS m3_n2650_n13200# m3_n7969_n2600# m3_7988_8000#
+ m3_2669_n7900# m3_n13288_n2600# m3_n2650_2700# m3_2669_2700# m3_n13288_n13200# m3_n7969_n13200#
+ m3_n13288_8000# m3_7988_2700# m3_n2650_n7900# m3_7988_n7900# m3_2669_n13200# m3_n7969_8000#
+ m3_n13288_2700# m3_n7969_n7900# m3_n13288_n7900# m3_2669_n2600# m3_n7969_2700# m3_7988_n13200#
+ c1_n13188_n13100# m3_7988_n2600# m3_n2650_n2600# m3_n2650_8000# m3_2669_8000#
X0 c1_n13188_n13100# m3_2669_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X1 c1_n13188_n13100# m3_n2650_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X2 c1_n13188_n13100# m3_2669_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X3 c1_n13188_n13100# m3_n13288_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X4 c1_n13188_n13100# m3_n7969_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X5 c1_n13188_n13100# m3_n13288_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X6 c1_n13188_n13100# m3_2669_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X7 c1_n13188_n13100# m3_7988_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X8 c1_n13188_n13100# m3_2669_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X9 c1_n13188_n13100# m3_7988_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X10 c1_n13188_n13100# m3_n7969_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X11 c1_n13188_n13100# m3_7988_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X12 c1_n13188_n13100# m3_n7969_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X13 c1_n13188_n13100# m3_7988_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X14 c1_n13188_n13100# m3_n13288_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X15 c1_n13188_n13100# m3_n7969_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X16 c1_n13188_n13100# m3_n2650_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X17 c1_n13188_n13100# m3_n2650_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X18 c1_n13188_n13100# m3_n2650_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X19 c1_n13188_n13100# m3_7988_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X20 c1_n13188_n13100# m3_n13288_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X21 c1_n13188_n13100# m3_n13288_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X22 c1_n13188_n13100# m3_n7969_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X23 c1_n13188_n13100# m3_n2650_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X24 c1_n13188_n13100# m3_2669_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
C0 m3_n7969_n13200# c1_n13188_n13100# 58.61fF
C1 c1_n13188_n13100# m3_n2650_n13200# 58.61fF
C2 c1_n13188_n13100# m3_n2650_8000# 58.61fF
C3 m3_7988_2700# c1_n13188_n13100# 61.01fF
C4 m3_n2650_2700# c1_n13188_n13100# 58.86fF
C5 m3_n2650_n13200# m3_2669_n13200# 2.73fF
C6 c1_n13188_n13100# m3_2669_8000# 58.61fF
C7 m3_n7969_2700# m3_n13288_2700# 2.73fF
C8 m3_7988_8000# c1_n13188_n13100# 60.75fF
C9 m3_n13288_n7900# m3_n13288_n13200# 3.28fF
C10 m3_n13288_8000# c1_n13188_n13100# 58.36fF
C11 m3_7988_n7900# c1_n13188_n13100# 61.01fF
C12 m3_n7969_8000# m3_n2650_8000# 2.73fF
C13 m3_n2650_n7900# m3_n2650_n13200# 3.28fF
C14 c1_n13188_n13100# m3_n7969_n7900# 58.86fF
C15 m3_n13288_n2600# m3_n13288_2700# 3.28fF
C16 m3_n13288_8000# m3_n7969_8000# 2.73fF
C17 m3_7988_n7900# m3_2669_n7900# 2.73fF
C18 m3_7988_2700# m3_2669_2700# 2.73fF
C19 m3_n7969_n7900# m3_n2650_n7900# 2.73fF
C20 m3_n7969_n2600# m3_n7969_n7900# 3.28fF
C21 m3_n2650_2700# m3_2669_2700# 2.73fF
C22 c1_n13188_n13100# m3_2669_n13200# 58.61fF
C23 m3_2669_8000# m3_2669_2700# 3.28fF
C24 m3_n13288_n7900# m3_n7969_n7900# 2.73fF
C25 c1_n13188_n13100# m3_n7969_8000# 58.61fF
C26 m3_n2650_2700# m3_n2650_n2600# 3.28fF
C27 c1_n13188_n13100# m3_2669_n7900# 58.86fF
C28 c1_n13188_n13100# m3_n2650_n7900# 58.86fF
C29 m3_n7969_n2600# c1_n13188_n13100# 58.86fF
C30 m3_2669_n7900# m3_2669_n13200# 3.28fF
C31 m3_n2650_2700# m3_n7969_2700# 2.73fF
C32 m3_n13288_n7900# c1_n13188_n13100# 58.61fF
C33 c1_n13188_n13100# m3_2669_n2600# 58.86fF
C34 m3_7988_n2600# m3_7988_2700# 3.39fF
C35 c1_n13188_n13100# m3_2669_2700# 58.86fF
C36 m3_n2650_n7900# m3_2669_n7900# 2.73fF
C37 m3_n13288_8000# m3_n13288_2700# 3.28fF
C38 m3_7988_n7900# m3_7988_n13200# 3.39fF
C39 m3_2669_n7900# m3_2669_n2600# 3.28fF
C40 m3_n2650_n2600# c1_n13188_n13100# 58.86fF
C41 m3_7988_n2600# m3_7988_n7900# 3.39fF
C42 m3_n7969_2700# c1_n13188_n13100# 58.86fF
C43 m3_n7969_n13200# m3_n13288_n13200# 2.73fF
C44 m3_7988_n13200# c1_n13188_n13100# 60.75fF
C45 c1_n13188_n13100# m3_n13288_2700# 58.61fF
C46 m3_2669_2700# m3_2669_n2600# 3.28fF
C47 m3_n2650_n2600# m3_n2650_n7900# 3.28fF
C48 m3_n13288_n2600# c1_n13188_n13100# 58.61fF
C49 m3_n7969_n13200# m3_n2650_n13200# 2.73fF
C50 m3_n7969_n2600# m3_n2650_n2600# 2.73fF
C51 m3_7988_n2600# c1_n13188_n13100# 61.01fF
C52 m3_7988_n13200# m3_2669_n13200# 2.73fF
C53 m3_n7969_2700# m3_n7969_8000# 3.28fF
C54 m3_n2650_n2600# m3_2669_n2600# 2.73fF
C55 m3_n7969_n2600# m3_n7969_2700# 3.28fF
C56 m3_n2650_2700# m3_n2650_8000# 3.28fF
C57 m3_2669_8000# m3_n2650_8000# 2.73fF
C58 m3_n7969_n2600# m3_n13288_n2600# 2.73fF
C59 m3_n7969_n13200# m3_n7969_n7900# 3.28fF
C60 m3_7988_2700# m3_7988_8000# 3.39fF
C61 m3_n13288_n7900# m3_n13288_n2600# 3.28fF
C62 m3_7988_n2600# m3_2669_n2600# 2.73fF
C63 m3_7988_8000# m3_2669_8000# 2.73fF
C64 c1_n13188_n13100# m3_n13288_n13200# 58.36fF
C65 c1_n13188_n13100# VSUBS 2.51fF
C66 m3_7988_n13200# VSUBS 12.57fF
C67 m3_2669_n13200# VSUBS 12.37fF
C68 m3_n2650_n13200# VSUBS 12.37fF
C69 m3_n7969_n13200# VSUBS 12.37fF
C70 m3_n13288_n13200# VSUBS 12.37fF
C71 m3_7988_n7900# VSUBS 12.57fF
C72 m3_2669_n7900# VSUBS 12.37fF
C73 m3_n2650_n7900# VSUBS 12.37fF
C74 m3_n7969_n7900# VSUBS 12.37fF
C75 m3_n13288_n7900# VSUBS 12.37fF
C76 m3_7988_n2600# VSUBS 12.57fF
C77 m3_2669_n2600# VSUBS 12.37fF
C78 m3_n2650_n2600# VSUBS 12.37fF
C79 m3_n7969_n2600# VSUBS 12.37fF
C80 m3_n13288_n2600# VSUBS 12.37fF
C81 m3_7988_2700# VSUBS 12.57fF
C82 m3_2669_2700# VSUBS 12.37fF
C83 m3_n2650_2700# VSUBS 12.37fF
C84 m3_n7969_2700# VSUBS 12.37fF
C85 m3_n13288_2700# VSUBS 12.37fF
C86 m3_7988_8000# VSUBS 12.57fF
C87 m3_2669_8000# VSUBS 12.37fF
C88 m3_n2650_8000# VSUBS 12.37fF
C89 m3_n7969_8000# VSUBS 12.37fF
C90 m3_n13288_8000# VSUBS 12.37fF
.ends

.subckt cap1_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_MACBVW_0 VSUBS out out out out out out out out out out
+ out out out out out out out out out out out in out out out out sky130_fd_pr__cap_mim_m3_1_MACBVW
C0 in out 2.17fF
C1 in VSUBS -10.03fF
C2 out VSUBS 62.40fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WHJTNJ VSUBS m3_n4309_50# m3_n4309_n4250# c1_n4209_n4150#
+ c1_110_n4150# m3_10_n4250#
X0 c1_n4209_n4150# m3_n4309_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 c1_110_n4150# m3_10_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2 c1_n4209_n4150# m3_n4309_50# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 c1_110_n4150# m3_10_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
C0 c1_n4209_n4150# c1_110_n4150# 1.32fF
C1 m3_n4309_n4250# m3_10_n4250# 1.75fF
C2 c1_n4209_n4150# m3_n4309_50# 38.10fF
C3 m3_n4309_50# m3_n4309_n4250# 2.63fF
C4 c1_n4209_n4150# m3_n4309_n4250# 38.10fF
C5 c1_110_n4150# m3_10_n4250# 81.11fF
C6 m3_n4309_50# m3_10_n4250# 1.75fF
C7 c1_110_n4150# VSUBS 0.12fF
C8 c1_n4209_n4150# VSUBS 0.12fF
C9 m3_n4309_n4250# VSUBS 8.68fF
C10 m3_10_n4250# VSUBS 17.92fF
C11 m3_n4309_50# VSUBS 8.68fF
.ends

.subckt cap3_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_WHJTNJ_0 VSUBS out out in in out sky130_fd_pr__cap_mim_m3_1_WHJTNJ
C0 in out 3.21fF
C1 in VSUBS -8.91fF
C2 out VSUBS 3.92fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_W3JTNJ VSUBS m3_n6469_n2100# c1_n6369_n6300# m3_2169_n6400#
+ m3_n2150_n6400# c1_2269_n6300# m3_n6469_2200# m3_n2150_n2100# c1_n2050_n6300# m3_n2150_2200#
+ m3_n6469_n6400#
X0 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2 c1_n2050_n6300# m3_n2150_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 c1_n6369_n6300# m3_n6469_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X4 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X5 c1_n6369_n6300# m3_n6469_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X6 c1_n2050_n6300# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X7 c1_n2050_n6300# m3_n2150_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X8 c1_n6369_n6300# m3_n6469_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
C0 m3_n2150_2200# m3_n6469_2200# 1.75fF
C1 c1_n6369_n6300# c1_n2050_n6300# 1.99fF
C2 m3_n2150_n6400# m3_n2150_n2100# 2.63fF
C3 m3_2169_n6400# m3_n2150_n6400# 1.75fF
C4 c1_n6369_n6300# m3_n6469_2200# 38.10fF
C5 m3_n2150_n2100# c1_n2050_n6300# 38.10fF
C6 m3_n2150_n6400# m3_n6469_n6400# 1.75fF
C7 m3_n2150_2200# m3_n2150_n2100# 2.63fF
C8 c1_2269_n6300# m3_2169_n6400# 121.67fF
C9 m3_n2150_2200# m3_2169_n6400# 1.75fF
C10 m3_n6469_n2100# m3_n6469_2200# 2.63fF
C11 m3_n6469_n2100# c1_n6369_n6300# 38.10fF
C12 m3_n2150_n6400# c1_n2050_n6300# 38.10fF
C13 c1_n6369_n6300# m3_n6469_n6400# 38.10fF
C14 m3_n6469_n2100# m3_n2150_n2100# 1.75fF
C15 m3_2169_n6400# m3_n2150_n2100# 1.75fF
C16 c1_2269_n6300# c1_n2050_n6300# 1.99fF
C17 m3_n2150_2200# c1_n2050_n6300# 38.10fF
C18 m3_n6469_n2100# m3_n6469_n6400# 2.63fF
C19 c1_2269_n6300# VSUBS 0.16fF
C20 c1_n2050_n6300# VSUBS 0.16fF
C21 c1_n6369_n6300# VSUBS 0.16fF
C22 m3_n2150_n6400# VSUBS 8.68fF
C23 m3_n6469_n6400# VSUBS 8.68fF
C24 m3_n2150_n2100# VSUBS 8.68fF
C25 m3_n6469_n2100# VSUBS 8.68fF
C26 m3_2169_n6400# VSUBS 26.86fF
C27 m3_n2150_2200# VSUBS 8.68fF
C28 m3_n6469_2200# VSUBS 8.68fF
.ends

.subckt cap2_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_W3JTNJ_0 VSUBS out in out out in out out in out out sky130_fd_pr__cap_mim_m3_1_W3JTNJ
C0 in out 8.08fF
C1 in VSUBS -16.59fF
C2 out VSUBS 13.00fF
.ends

.subckt sky130_fd_pr__nfet_01v8_U2JGXT w_n226_n510# a_n118_n388# a_n88_n300# a_30_n300#
X0 a_30_n300# a_n118_n388# a_n88_n300# w_n226_n510# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
C0 a_n88_n300# a_n118_n388# 0.11fF
C1 a_n88_n300# a_30_n300# 0.61fF
C2 a_30_n300# w_n226_n510# 0.40fF
C3 a_n88_n300# w_n226_n510# 0.40fF
C4 a_n118_n388# w_n226_n510# 0.28fF
.ends

.subckt sky130_fd_pr__res_high_po_5p73_X44RQA a_n573_2292# w_n739_n2890# a_n573_n2724#
X0 a_n573_n2724# a_n573_2292# w_n739_n2890# sky130_fd_pr__res_high_po_5p73 l=2.292e+07u
C0 a_n573_n2724# w_n739_n2890# 1.98fF
C1 a_n573_2292# w_n739_n2890# 1.98fF
.ends

.subckt res_loop_filter vss out in
Xsky130_fd_pr__res_high_po_5p73_X44RQA_0 in vss out sky130_fd_pr__res_high_po_5p73_X44RQA
C0 out vss 3.87fF
C1 in vss 3.02fF
.ends

.subckt loop_filter_v2 vc_pex D0_cap in vss cap3_loop_filter_0/in
Xcap1_loop_filter_0 vss vc_pex vss cap1_loop_filter
Xcap3_loop_filter_0 vss cap3_loop_filter_0/in vss cap3_loop_filter
Xcap2_loop_filter_0 vss in vss cap2_loop_filter
Xsky130_fd_pr__nfet_01v8_U2JGXT_0 vss D0_cap in cap3_loop_filter_0/in sky130_fd_pr__nfet_01v8_U2JGXT
Xres_loop_filter_0 vss res_loop_filter_2/out in res_loop_filter
Xres_loop_filter_1 vss res_loop_filter_2/out vc_pex res_loop_filter
Xres_loop_filter_2 vss res_loop_filter_2/out vc_pex res_loop_filter
C0 cap3_loop_filter_0/in in 0.79fF
C1 in D0_cap 0.07fF
C2 vc_pex in 0.18fF
C3 vc_pex vss -38.13fF
C4 res_loop_filter_2/out vss 8.49fF
C5 D0_cap vss 0.04fF
C6 in vss -18.54fF
C7 cap3_loop_filter_0/in vss -3.74fF
.ends

.subckt sky130_fd_pr__pfet_01v8_58ZKDE VSUBS a_n257_n777# a_n129_n600# a_n221_n600#
+ w_n257_n702#
X0 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X1 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X2 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X3 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
C0 a_n257_n777# a_n221_n600# 0.25fF
C1 a_n221_n600# a_n129_n600# 7.87fF
C2 a_n257_n777# a_n129_n600# 0.29fF
C3 a_n129_n600# VSUBS 0.10fF
C4 a_n221_n600# VSUBS 0.25fF
C5 a_n257_n777# VSUBS 1.05fF
C6 w_n257_n702# VSUBS 2.16fF
.ends

.subckt sky130_fd_pr__nfet_01v8_T69Y3A a_n129_n300# a_n221_n300# w_n257_n327# a_n257_n404#
X0 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
C0 a_n221_n300# a_n129_n300# 4.05fF
C1 a_n257_n404# a_n129_n300# 0.30fF
C2 a_n257_n404# a_n221_n300# 0.21fF
C3 a_n129_n300# w_n257_n327# 0.11fF
C4 a_n221_n300# w_n257_n327# 0.25fF
C5 a_n257_n404# w_n257_n327# 1.11fF
.ends

.subckt buffer_salida a_678_n100# a_3996_n100# out vdd in vss
Xsky130_fd_pr__pfet_01v8_58ZKDE_1 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_2 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_3 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_0 a_678_n100# vss vss in sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_1 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_4 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_5 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_2 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_3 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_6 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_70 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_4 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_7 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_8 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_71 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_60 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_5 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_72 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_61 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_50 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_6 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_9 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_62 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_51 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_7 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_40 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_8 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_63 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_52 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_30 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_41 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_64 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_53 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_9 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_20 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_31 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_42 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_65 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_54 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_10 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_21 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_32 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_43 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_66 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_55 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_11 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_22 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_33 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_44 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_67 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_56 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_12 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_23 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_34 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_45 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_68 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_57 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_13 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_24 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_35 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_46 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_69 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_58 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_14 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_25 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_36 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_47 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_59 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_48 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_15 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_26 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_37 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_49 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_16 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_27 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_38 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_70 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_17 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_28 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_39 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_71 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_60 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_18 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_29 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_72 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_61 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_50 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_62 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_51 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_19 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_40 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_63 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_52 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_30 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_41 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_64 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_53 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_20 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_31 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_42 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_65 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_54 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_10 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_21 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_32 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_43 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_66 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_55 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_11 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_22 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_33 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_44 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_67 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_56 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_12 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_23 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_34 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_45 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_68 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_57 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_46 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_13 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_24 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_35 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_69 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_58 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_14 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_25 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_36 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_47 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_59 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_15 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_26 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_37 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_48 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_49 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_16 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_27 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_38 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_17 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_28 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_39 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_18 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_29 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_19 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_0 vss in a_678_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
C0 vdd a_678_n100# 0.08fF
C1 a_678_n100# a_3996_n100# 6.52fF
C2 vdd a_3996_n100# 3.68fF
C3 vdd out 47.17fF
C4 in a_678_n100# 0.81fF
C5 vdd in 0.02fF
C6 out a_3996_n100# 55.19fF
C7 vdd vss 20.93fF
C8 out vss 35.17fF
C9 a_3996_n100# vss 49.53fF
C10 a_678_n100# vss 13.08fF
C11 in vss 0.87fF
.ends

.subckt trans_gate_mux2to8 in vss out en_pos en_neg vdd
Xsky130_fd_pr__pfet_01v8_4798MH_0 vss en_neg in out out vdd en_neg en_neg in sky130_fd_pr__pfet_01v8_4798MH
Xsky130_fd_pr__nfet_01v8_BHR94T_0 en_pos vss en_pos in out out en_pos in sky130_fd_pr__nfet_01v8_BHR94T
C0 in vdd 0.05fF
C1 out en_neg 0.07fF
C2 vdd en_neg 0.01fF
C3 out en_pos 0.27fF
C4 in en_neg 0.28fF
C5 in en_pos 0.07fF
C6 out vdd 0.68fF
C7 en_pos en_neg 0.04fF
C8 out in 0.36fF
C9 vdd vss 2.75fF
C10 en_pos vss 0.30fF
C11 in vss 1.53fF
C12 out vss 0.88fF
C13 en_neg vss 0.31fF
.ends

.subckt mux2to1 vss select_0_neg in_a out_a_0 out_a_1 select_0 vdd
Xtrans_gate_mux2to8_0 in_a vss out_a_0 select_0_neg select_0 vdd trans_gate_mux2to8
Xtrans_gate_mux2to8_1 in_a vss out_a_1 select_0 select_0_neg vdd trans_gate_mux2to8
C0 vdd out_a_1 0.09fF
C1 select_0 in_a 0.31fF
C2 select_0 select_0_neg 0.17fF
C3 out_a_0 vdd 0.09fF
C4 in_a select_0_neg 0.11fF
C5 select_0 vdd 0.04fF
C6 in_a vdd 0.14fF
C7 select_0 out_a_1 0.14fF
C8 in_a out_a_1 0.08fF
C9 in_a out_a_0 0.08fF
C10 select_0_neg out_a_0 0.05fF
C11 out_a_1 vss 1.03fF
C12 vdd vss 6.09fF
C13 select_0_neg vss 1.12fF
C14 in_a vss 2.43fF
C15 out_a_0 vss 1.03fF
C16 select_0 vss 1.03fF
.ends

.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X a_194_125# a_355_368# a_455_87#
+ a_158_392#
X0 X B a_455_87# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 X a_194_125# a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_194_125# B a_158_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_158_392# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_355_368# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_194_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 a_455_87# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND B a_194_125# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X9 VGND a_194_125# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
C0 a_194_125# A 0.18fF
C1 A VPWR 0.15fF
C2 a_158_392# a_194_125# 0.06fF
C3 a_194_125# VPWR 0.33fF
C4 a_194_125# X 0.29fF
C5 X VPWR 0.07fF
C6 A VGND 0.31fF
C7 a_194_125# VGND 0.25fF
C8 VGND VPWR 0.01fF
C9 X VGND 0.28fF
C10 A B 0.28fF
C11 VPWR VPB 0.06fF
C12 a_194_125# B 0.57fF
C13 VPWR B 0.09fF
C14 A a_355_368# 0.02fF
C15 a_194_125# a_355_368# 0.51fF
C16 VPWR a_355_368# 0.37fF
C17 X B 0.13fF
C18 VGND B 0.10fF
C19 X a_355_368# 0.17fF
C20 B a_355_368# 0.08fF
C21 VGND VNB 0.78fF
C22 X VNB 0.21fF
C23 VPWR VNB 0.78fF
C24 B VNB 0.56fF
C25 A VNB 0.70fF
C26 VPB VNB 0.77fF
C27 a_355_368# VNB 0.08fF
C28 a_194_125# VNB 0.40fF
.ends

.subckt sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X a_143_136# a_56_136#
X0 VGND B a_143_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 X a_56_136# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VPWR B a_56_136# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_143_136# A a_56_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_56_136# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 X a_56_136# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
C0 VPWR A 0.07fF
C1 A a_56_136# 0.17fF
C2 VPWR a_56_136# 0.57fF
C3 VGND B 0.03fF
C4 VGND X 0.15fF
C5 VPWR VPB 0.04fF
C6 A B 0.08fF
C7 VPWR B 0.02fF
C8 X VPWR 0.20fF
C9 a_56_136# B 0.30fF
C10 X a_56_136# 0.26fF
C11 VGND A 0.21fF
C12 VGND a_56_136# 0.06fF
C13 X B 0.02fF
C14 VGND VNB 0.50fF
C15 X VNB 0.23fF
C16 VPWR VNB 0.50fF
C17 B VNB 0.24fF
C18 A VNB 0.36fF
C19 VPB VNB 0.48fF
C20 a_56_136# VNB 0.38fF
.ends

.subckt sky130_fd_sc_hs__or2_1 A B VGND VNB VPB VPWR X a_152_368# a_63_368#
X0 VPWR A a_152_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_152_368# B a_63_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 X a_63_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 X a_63_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_63_368# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X5 VGND A a_63_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
C0 a_63_368# A 0.28fF
C1 X A 0.02fF
C2 B A 0.10fF
C3 VPWR a_63_368# 0.29fF
C4 VPWR X 0.18fF
C5 VPWR B 0.01fF
C6 X a_63_368# 0.33fF
C7 a_63_368# B 0.14fF
C8 VPWR VPB 0.04fF
C9 a_63_368# VGND 0.27fF
C10 X VGND 0.16fF
C11 B VGND 0.11fF
C12 VPWR A 0.05fF
C13 a_63_368# a_152_368# 0.03fF
C14 VGND VNB 0.53fF
C15 X VNB 0.24fF
C16 A VNB 0.21fF
C17 B VNB 0.31fF
C18 VPWR VNB 0.46fF
C19 VPB VNB 0.48fF
C20 a_63_368# VNB 0.37fF
.ends

.subckt div_by_5 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in nCLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_0/latch_diff_1/nD vss vdd DFlipFlop_2/latch_diff_0/nD Q0 Q1 CLK DFlipFlop_0/Q
+ DFlipFlop_2/latch_diff_1/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out sky130_fd_sc_hs__and2_1_0/a_56_136#
+ nQ0 DFlipFlop_3/latch_diff_0/D DFlipFlop_3/latch_diff_1/nD DFlipFlop_1/latch_diff_1/nD
+ DFlipFlop_1/latch_diff_0/nD DFlipFlop_1/latch_diff_0/D DFlipFlop_2/latch_diff_0/m1_657_280#
+ CLK_5 Q1_shift nQ2 DFlipFlop_2/D DFlipFlop_2/latch_diff_1/nD DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_1/latch_diff_1/D DFlipFlop_1/D DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_0/latch_diff_0/nD sky130_fd_sc_hs__xor2_1_0/a_355_368# DFlipFlop_0/D DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_0/latch_diff_1/D DFlipFlop_2/nQ DFlipFlop_3/latch_diff_0/nD DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_2/latch_diff_0/D DFlipFlop_0/latch_diff_0/D sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ DFlipFlop_3/latch_diff_1/D sky130_fd_sc_hs__or2_1_0/a_63_368# DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ sky130_fd_sc_hs__and2_1_1/a_143_136# sky130_fd_sc_hs__or2_1_0/a_152_368# sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ sky130_fd_sc_hs__and2_1_1/a_56_136# DFlipFlop_3/nQ sky130_fd_sc_hs__and2_1_0/a_143_136#
Xsky130_fd_sc_hs__xor2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_2/D sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ sky130_fd_sc_hs__xor2_1_0/a_355_368# sky130_fd_sc_hs__xor2_1_0/a_455_87# sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ sky130_fd_sc_hs__xor2_1
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vss vdd DFlipFlop_0/latch_diff_1/D
+ DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in nQ2 nCLK DFlipFlop_0/latch_diff_0/nD
+ DFlipFlop_0/Q DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/latch_diff_1/m1_657_280# DFlipFlop_0/D
+ DFlipFlop_0/latch_diff_0/D CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_1 DFlipFlop_1/latch_diff_0/m1_657_280# vss vdd DFlipFlop_1/latch_diff_1/D
+ DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in nQ0 nCLK DFlipFlop_1/latch_diff_0/nD
+ Q0 DFlipFlop_1/latch_diff_1/nD DFlipFlop_1/latch_diff_1/m1_657_280# DFlipFlop_1/D
+ DFlipFlop_1/latch_diff_0/D CLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_2 DFlipFlop_2/latch_diff_0/m1_657_280# vss vdd DFlipFlop_2/latch_diff_1/D
+ DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_2/nQ nCLK DFlipFlop_2/latch_diff_0/nD
+ Q1 DFlipFlop_2/latch_diff_1/nD DFlipFlop_2/latch_diff_1/m1_657_280# DFlipFlop_2/D
+ DFlipFlop_2/latch_diff_0/D CLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_3 DFlipFlop_3/latch_diff_0/m1_657_280# vss vdd DFlipFlop_3/latch_diff_1/D
+ DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_3/nQ CLK DFlipFlop_3/latch_diff_0/nD
+ Q1_shift DFlipFlop_3/latch_diff_1/nD DFlipFlop_3/latch_diff_1/m1_657_280# Q1 DFlipFlop_3/latch_diff_0/D
+ nCLK DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop
Xsky130_fd_sc_hs__and2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_0/D sky130_fd_sc_hs__and2_1_0/a_143_136#
+ sky130_fd_sc_hs__and2_1_0/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__and2_1_1 nQ2 nQ0 vss vss vdd vdd DFlipFlop_1/D sky130_fd_sc_hs__and2_1_1/a_143_136#
+ sky130_fd_sc_hs__and2_1_1/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__or2_1_0 Q1 Q1_shift vss vss vdd vdd CLK_5 sky130_fd_sc_hs__or2_1_0/a_152_368#
+ sky130_fd_sc_hs__or2_1_0/a_63_368# sky130_fd_sc_hs__or2_1
C0 vdd nCLK 0.34fF
C1 sky130_fd_sc_hs__or2_1_0/a_152_368# Q1_shift -0.04fF
C2 DFlipFlop_2/nQ nCLK 0.09fF
C3 DFlipFlop_1/D Q1 0.03fF
C4 DFlipFlop_1/latch_diff_1/D Q1 -0.10fF
C5 DFlipFlop_3/latch_diff_0/m1_657_280# nCLK 0.27fF
C6 DFlipFlop_2/latch_diff_1/m1_657_280# nCLK 0.28fF
C7 CLK vdd 0.41fF
C8 CLK DFlipFlop_1/latch_diff_0/m1_657_280# 0.28fF
C9 DFlipFlop_2/latch_diff_0/D Q1 0.42fF
C10 CLK DFlipFlop_2/nQ 0.13fF
C11 DFlipFlop_2/latch_diff_1/D Q1 0.23fF
C12 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in nCLK 0.14fF
C13 sky130_fd_sc_hs__or2_1_0/a_63_368# Q1 0.10fF
C14 DFlipFlop_2/D sky130_fd_sc_hs__xor2_1_0/a_194_125# 0.08fF
C15 DFlipFlop_0/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.02fF
C16 sky130_fd_sc_hs__xor2_1_0/a_455_87# nCLK 0.02fF
C17 Q1 nCLK -0.01fF
C18 CLK DFlipFlop_2/latch_diff_0/m1_657_280# 0.28fF
C19 DFlipFlop_1/latch_diff_0/D Q1 0.18fF
C20 vdd DFlipFlop_0/D 0.19fF
C21 sky130_fd_sc_hs__xor2_1_0/a_194_125# Q0 0.26fF
C22 DFlipFlop_1/latch_diff_1/nD nCLK 0.16fF
C23 DFlipFlop_2/D Q0 0.25fF
C24 DFlipFlop_0/Q Q0 0.21fF
C25 DFlipFlop_3/latch_diff_1/nD nCLK 0.09fF
C26 nQ0 DFlipFlop_1/D 0.12fF
C27 DFlipFlop_3/nQ nCLK 0.02fF
C28 nQ0 DFlipFlop_1/latch_diff_1/D 0.91fF
C29 nQ2 DFlipFlop_0/Q 0.09fF
C30 CLK Q1 -0.10fF
C31 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vdd 0.03fF
C32 nQ0 DFlipFlop_1/latch_diff_1/m1_657_280# 0.21fF
C33 DFlipFlop_1/latch_diff_1/nD CLK 0.09fF
C34 nQ2 Q0 0.23fF
C35 vdd Q1_shift 0.10fF
C36 sky130_fd_sc_hs__and2_1_1/a_143_136# CLK 0.03fF
C37 DFlipFlop_3/latch_diff_1/nD CLK 0.16fF
C38 DFlipFlop_0/latch_diff_1/m1_657_280# nCLK 0.28fF
C39 CLK DFlipFlop_3/nQ 0.01fF
C40 DFlipFlop_3/latch_diff_1/D Q1 0.79fF
C41 Q1 DFlipFlop_0/D 0.13fF
C42 DFlipFlop_0/latch_diff_0/D Q0 0.42fF
C43 CLK DFlipFlop_3/latch_diff_0/D 0.11fF
C44 DFlipFlop_0/latch_diff_1/D CLK 0.03fF
C45 nQ2 sky130_fd_sc_hs__and2_1_1/a_56_136# 0.01fF
C46 CLK DFlipFlop_3/latch_diff_1/m1_657_280# 0.27fF
C47 nQ0 nCLK 0.09fF
C48 DFlipFlop_1/latch_diff_0/D nQ0 0.09fF
C49 sky130_fd_sc_hs__and2_1_0/a_56_136# DFlipFlop_0/D 0.04fF
C50 Q1 DFlipFlop_3/latch_diff_0/nD 0.08fF
C51 sky130_fd_sc_hs__xor2_1_0/a_194_125# vdd 0.03fF
C52 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in Q1 0.20fF
C53 CLK_5 sky130_fd_sc_hs__or2_1_0/a_63_368# 0.06fF
C54 DFlipFlop_0/latch_diff_1/nD nCLK 0.05fF
C55 DFlipFlop_2/D vdd 0.07fF
C56 Q1 DFlipFlop_2/latch_diff_1/nD 0.21fF
C57 Q1 Q1_shift 0.36fF
C58 nQ0 CLK 0.19fF
C59 vdd DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C60 Q0 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.33fF
C61 DFlipFlop_1/D nCLK 0.14fF
C62 DFlipFlop_1/latch_diff_1/D nCLK 0.08fF
C63 vdd Q0 5.33fF
C64 nQ2 vdd 0.04fF
C65 DFlipFlop_0/latch_diff_1/nD CLK 0.02fF
C66 DFlipFlop_1/latch_diff_1/m1_657_280# nCLK 0.28fF
C67 DFlipFlop_3/nQ Q1_shift 0.04fF
C68 DFlipFlop_2/latch_diff_0/D nCLK 0.11fF
C69 DFlipFlop_2/latch_diff_1/D nCLK 0.08fF
C70 DFlipFlop_1/D CLK 0.21fF
C71 DFlipFlop_1/latch_diff_1/D CLK 0.14fF
C72 vdd sky130_fd_sc_hs__and2_1_1/a_56_136# 0.04fF
C73 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vdd 0.02fF
C74 DFlipFlop_2/D sky130_fd_sc_hs__xor2_1_0/a_455_87# 0.08fF
C75 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in Q0 0.42fF
C76 DFlipFlop_2/D Q1 0.10fF
C77 DFlipFlop_0/Q Q1 0.13fF
C78 sky130_fd_sc_hs__and2_1_0/a_143_136# Q0 0.03fF
C79 Q1 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out 0.15fF
C80 CLK DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in 0.03fF
C81 DFlipFlop_1/latch_diff_0/D nCLK 0.11fF
C82 DFlipFlop_2/latch_diff_1/D CLK 0.14fF
C83 Q1 Q0 9.65fF
C84 nQ2 Q1 0.07fF
C85 vdd DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.02fF
C86 DFlipFlop_1/latch_diff_1/nD Q0 0.21fF
C87 sky130_fd_sc_hs__and2_1_0/a_56_136# Q0 0.17fF
C88 DFlipFlop_0/latch_diff_0/D Q1 0.15fF
C89 nQ2 sky130_fd_sc_hs__and2_1_1/a_143_136# 0.01fF
C90 DFlipFlop_2/nQ vdd 0.02fF
C91 DFlipFlop_0/latch_diff_1/D Q0 0.23fF
C92 sky130_fd_sc_hs__xor2_1_0/a_355_368# Q0 0.03fF
C93 DFlipFlop_3/latch_diff_1/D nCLK 0.14fF
C94 CLK DFlipFlop_0/latch_diff_0/m1_657_280# 0.28fF
C95 nQ2 DFlipFlop_0/latch_diff_1/m1_657_280# 0.05fF
C96 nCLK DFlipFlop_3/latch_diff_0/nD 0.08fF
C97 Q1 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.09fF
C98 sky130_fd_sc_hs__or2_1_0/a_63_368# Q1_shift -0.27fF
C99 CLK DFlipFlop_3/latch_diff_1/D 0.08fF
C100 nQ0 Q0 0.33fF
C101 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in nCLK -0.33fF
C102 vdd Q1 9.49fF
C103 nQ2 nQ0 0.03fF
C104 DFlipFlop_2/nQ Q1 0.31fF
C105 nCLK DFlipFlop_2/latch_diff_1/nD 0.16fF
C106 CLK DFlipFlop_2/latch_diff_0/nD 0.08fF
C107 DFlipFlop_3/latch_diff_0/m1_657_280# Q1 0.28fF
C108 DFlipFlop_1/latch_diff_0/nD nQ0 0.08fF
C109 DFlipFlop_0/latch_diff_1/nD Q0 0.21fF
C110 nQ0 sky130_fd_sc_hs__and2_1_1/a_56_136# 0.01fF
C111 sky130_fd_sc_hs__and2_1_0/a_56_136# vdd 0.02fF
C112 vdd DFlipFlop_3/nQ 0.02fF
C113 DFlipFlop_2/latch_diff_1/m1_657_280# Q1 0.03fF
C114 DFlipFlop_2/D DFlipFlop_1/latch_diff_1/m1_657_280# 0.04fF
C115 DFlipFlop_1/D Q0 0.07fF
C116 DFlipFlop_1/latch_diff_1/D Q0 0.06fF
C117 Q1 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in 0.21fF
C118 CLK DFlipFlop_2/latch_diff_1/nD 0.09fF
C119 vdd sky130_fd_sc_hs__xor2_1_0/a_355_368# 0.03fF
C120 sky130_fd_sc_hs__and2_1_0/a_143_136# Q1 0.02fF
C121 DFlipFlop_1/latch_diff_1/m1_657_280# Q0 0.01fF
C122 sky130_fd_sc_hs__xor2_1_0/a_194_125# nCLK 0.11fF
C123 DFlipFlop_1/D DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C124 DFlipFlop_1/D sky130_fd_sc_hs__and2_1_1/a_56_136# 0.04fF
C125 DFlipFlop_2/D nCLK 0.41fF
C126 DFlipFlop_0/Q nCLK 0.11fF
C127 DFlipFlop_1/latch_diff_1/nD Q1 0.10fF
C128 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out nCLK 0.05fF
C129 nQ0 vdd 0.11fF
C130 sky130_fd_sc_hs__and2_1_0/a_56_136# Q1 0.14fF
C131 nQ0 DFlipFlop_1/latch_diff_0/m1_657_280# 0.25fF
C132 DFlipFlop_3/latch_diff_1/nD Q1 1.24fF
C133 Q1 DFlipFlop_3/nQ 0.10fF
C134 nCLK Q0 0.20fF
C135 DFlipFlop_1/latch_diff_0/D Q0 0.42fF
C136 nQ2 nCLK 0.10fF
C137 DFlipFlop_2/D CLK 0.14fF
C138 CLK DFlipFlop_0/Q 0.08fF
C139 Q1 DFlipFlop_3/latch_diff_0/D 0.09fF
C140 DFlipFlop_0/latch_diff_1/D Q1 0.06fF
C141 Q1 DFlipFlop_3/latch_diff_1/m1_657_280# 0.28fF
C142 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out CLK -0.31fF
C143 CLK_5 vdd 0.15fF
C144 CLK Q0 0.08fF
C145 DFlipFlop_1/D vdd 0.25fF
C146 nQ2 CLK 0.17fF
C147 nQ0 Q1 0.06fF
C148 DFlipFlop_1/latch_diff_0/nD CLK 0.08fF
C149 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vdd 0.03fF
C150 CLK sky130_fd_sc_hs__and2_1_1/a_56_136# 0.06fF
C151 CLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out 0.15fF
C152 sky130_fd_sc_hs__or2_1_0/a_63_368# vdd 0.02fF
C153 DFlipFlop_0/D Q0 0.39fF
C154 DFlipFlop_1/latch_diff_1/nD nQ0 0.88fF
C155 sky130_fd_sc_hs__and2_1_1/a_143_136# nQ0 0.04fF
C156 DFlipFlop_0/latch_diff_1/nD Q1 0.10fF
C157 CLK_5 vss -0.18fF
C158 sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.38fF
C159 sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.41fF
C160 sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C161 Q1_shift vss -0.29fF
C162 DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.64fF
C163 DFlipFlop_3/nQ vss 0.52fF
C164 DFlipFlop_3/latch_diff_1/D vss -1.73fF
C165 DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C166 DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C167 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.94fF
C168 DFlipFlop_3/latch_diff_0/D vss 0.96fF
C169 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.85fF
C170 DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C171 Q1 vss 8.55fF
C172 DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.72fF
C173 DFlipFlop_2/nQ vss 0.50fF
C174 DFlipFlop_2/latch_diff_1/D vss -1.72fF
C175 DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C176 DFlipFlop_2/latch_diff_1/nD vss 0.58fF
C177 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.89fF
C178 DFlipFlop_2/latch_diff_0/D vss 0.96fF
C179 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C180 DFlipFlop_2/D vss 5.34fF
C181 DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C182 Q0 vss 0.53fF
C183 DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.62fF
C184 nQ0 vss 3.42fF
C185 DFlipFlop_1/latch_diff_1/D vss -1.73fF
C186 DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C187 DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C188 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C189 DFlipFlop_1/latch_diff_0/D vss 0.96fF
C190 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.78fF
C191 DFlipFlop_1/D vss 3.72fF
C192 DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C193 DFlipFlop_0/Q vss -0.94fF
C194 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.61fF
C195 nCLK vss 0.96fF
C196 nQ2 vss 2.05fF
C197 DFlipFlop_0/latch_diff_1/D vss -1.73fF
C198 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C199 CLK vss 0.20fF
C200 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C201 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.88fF
C202 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C203 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C204 DFlipFlop_0/D vss 4.04fF
C205 vdd vss 146.76fF
C206 DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C207 sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C208 sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.42fF
.ends

.subckt mux2to4 vss out_b_1 vdd select_0 select_0_neg in_a out_a_0 out_a_1 out_b_0
+ in_b
Xtrans_gate_mux2to8_0 in_a vss out_a_0 select_0_neg select_0 vdd trans_gate_mux2to8
Xtrans_gate_mux2to8_1 in_a vss out_a_1 select_0 select_0_neg vdd trans_gate_mux2to8
Xtrans_gate_mux2to8_2 in_b vss out_b_0 select_0_neg select_0 vdd trans_gate_mux2to8
Xtrans_gate_mux2to8_3 in_b vss out_b_1 select_0 select_0_neg vdd trans_gate_mux2to8
C0 in_b select_0_neg 0.10fF
C1 out_b_0 out_a_1 0.88fF
C2 select_0_neg out_a_0 0.05fF
C3 in_b vdd 0.17fF
C4 select_0_neg select_0 0.49fF
C5 vdd out_a_0 0.09fF
C6 out_b_0 in_a 0.11fF
C7 in_a out_a_1 0.08fF
C8 vdd select_0 0.08fF
C9 select_0_neg vdd 0.08fF
C10 out_b_0 in_b 0.08fF
C11 in_b out_a_1 0.08fF
C12 in_b out_b_1 0.08fF
C13 out_b_0 select_0 0.03fF
C14 out_a_1 select_0 0.18fF
C15 out_b_0 select_0_neg -0.13fF
C16 select_0_neg out_a_1 0.12fF
C17 in_a out_a_0 0.08fF
C18 select_0 out_b_1 0.14fF
C19 in_a select_0 0.31fF
C20 out_b_0 vdd 0.15fF
C21 vdd out_a_1 0.16fF
C22 in_a select_0_neg 0.22fF
C23 vdd out_b_1 0.09fF
C24 in_a vdd 0.17fF
C25 in_b select_0 0.24fF
C26 out_b_1 vss 1.03fF
C27 in_b vss 2.46fF
C28 out_b_0 vss 0.84fF
C29 out_a_1 vss 0.32fF
C30 vdd vss 12.14fF
C31 select_0_neg vss 2.57fF
C32 in_a vss 2.46fF
C33 out_a_0 vss 1.03fF
C34 select_0 vss 2.24fF
.ends

.subckt sky130_fd_sc_hs__mux2_1 A0 A1 S VGND VNB VPB VPWR X a_304_74# a_443_74# a_524_368#
+ a_27_112#
X0 VPWR S a_27_112# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND a_27_112# a_443_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 X a_304_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VPWR a_27_112# a_524_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_304_74# A1 a_226_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 X a_304_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 a_223_368# S VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_304_74# A0 a_223_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_443_74# A0 a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_524_368# A1 a_304_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_226_74# S VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 VGND S a_27_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
C0 a_27_112# A0 0.07fF
C1 VPWR VGND 0.02fF
C2 VPWR A1 0.01fF
C3 a_223_368# a_304_74# 0.05fF
C4 VPWR a_304_74# 0.13fF
C5 a_443_74# A1 0.07fF
C6 VGND S 0.07fF
C7 S A1 0.10fF
C8 VGND A0 0.02fF
C9 A1 A0 0.31fF
C10 a_443_74# a_304_74# 0.12fF
C11 X a_27_112# 0.08fF
C12 VGND a_27_112# 0.18fF
C13 a_27_112# A1 0.18fF
C14 S a_304_74# 0.18fF
C15 A0 a_304_74# 0.23fF
C16 a_524_368# a_27_112# 0.06fF
C17 a_27_112# a_304_74# 0.58fF
C18 VPWR VPB 0.06fF
C19 VPWR S 0.05fF
C20 VGND X 0.11fF
C21 X A1 0.02fF
C22 VGND A1 0.09fF
C23 a_27_112# a_223_368# 0.09fF
C24 VPWR a_27_112# 0.99fF
C25 X a_304_74# 0.29fF
C26 a_226_74# a_304_74# 0.08fF
C27 VGND a_304_74# 0.58fF
C28 A1 a_304_74# 0.69fF
C29 S A0 0.04fF
C30 VPWR X 0.28fF
C31 a_27_112# VPB 0.01fF
C32 S a_27_112# 0.22fF
C33 VGND VNB 0.88fF
C34 X VNB 0.25fF
C35 VPWR VNB 0.89fF
C36 A1 VNB 0.37fF
C37 A0 VNB 0.23fF
C38 S VNB 0.34fF
C39 VPB VNB 0.87fF
C40 a_304_74# VNB 0.36fF
C41 a_27_112# VNB 0.65fF
.ends

.subckt prescaler_23 nCLK vss DFlipFlop_0/latch_diff_1/nD nCLK_23 DFlipFlop_2/latch_diff_0/nD
+ vdd DFlipFlop_2/latch_diff_1/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ CLK_23 DFlipFlop_2/latch_diff_0/m1_657_280# CLK DFlipFlop_2/latch_diff_1/nD DFlipFlop_0/latch_diff_0/nD
+ DFlipFlop_2/latch_diff_1/m1_657_280# DFlipFlop_0/latch_diff_1/D DFlipFlop_2/latch_diff_0/D
+ MC DFlipFlop_0/latch_diff_0/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in Q2
Xsky130_fd_sc_hs__mux2_1_0 sky130_fd_sc_hs__or2_1_1/X nCLK_23 MC vss vss vdd vdd CLK_23
+ sky130_fd_sc_hs__mux2_1_0/a_304_74# sky130_fd_sc_hs__mux2_1_0/a_443_74# sky130_fd_sc_hs__mux2_1_0/a_524_368#
+ sky130_fd_sc_hs__mux2_1_0/a_27_112# sky130_fd_sc_hs__mux2_1
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vss vdd DFlipFlop_0/latch_diff_1/D
+ DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_0/nQ nCLK DFlipFlop_0/latch_diff_0/nD
+ Q1 DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/latch_diff_1/m1_657_280# nCLK_23 DFlipFlop_0/latch_diff_0/D
+ CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop
XDFlipFlop_2 DFlipFlop_2/latch_diff_0/m1_657_280# vss vdd DFlipFlop_2/latch_diff_1/D
+ DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_2/nQ CLK DFlipFlop_2/latch_diff_0/nD
+ Q2_d DFlipFlop_2/latch_diff_1/nD DFlipFlop_2/latch_diff_1/m1_657_280# Q2 DFlipFlop_2/latch_diff_0/D
+ nCLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop
XDFlipFlop_1 DFlipFlop_1/latch_diff_0/m1_657_280# vss vdd DFlipFlop_1/latch_diff_1/D
+ DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in nCLK_23 nCLK DFlipFlop_1/latch_diff_0/nD
+ Q2 DFlipFlop_1/latch_diff_1/nD DFlipFlop_1/latch_diff_1/m1_657_280# DFlipFlop_1/D
+ DFlipFlop_1/latch_diff_0/D CLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
Xsky130_fd_sc_hs__and2_1_0 nCLK_23 sky130_fd_sc_hs__or2_1_0/X vss vss vdd vdd DFlipFlop_1/D
+ sky130_fd_sc_hs__and2_1_0/a_143_136# sky130_fd_sc_hs__and2_1_0/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__or2_1_0 Q1 MC vss vss vdd vdd sky130_fd_sc_hs__or2_1_0/X sky130_fd_sc_hs__or2_1_0/a_152_368#
+ sky130_fd_sc_hs__or2_1_0/a_63_368# sky130_fd_sc_hs__or2_1
Xsky130_fd_sc_hs__or2_1_1 Q2 Q2_d vss vss vdd vdd sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__or2_1_1/a_152_368#
+ sky130_fd_sc_hs__or2_1_1/a_63_368# sky130_fd_sc_hs__or2_1
C0 CLK DFlipFlop_1/latch_diff_1/nD 0.11fF
C1 nCLK DFlipFlop_2/nQ 0.02fF
C2 DFlipFlop_2/latch_diff_1/nD CLK 0.19fF
C3 sky130_fd_sc_hs__or2_1_0/X sky130_fd_sc_hs__and2_1_0/a_56_136# 0.07fF
C4 nCLK_23 DFlipFlop_0/latch_diff_1/nD 0.02fF
C5 MC Q1 0.29fF
C6 DFlipFlop_0/nQ Q1 -0.02fF
C7 sky130_fd_sc_hs__or2_1_0/X vdd 0.03fF
C8 CLK Q1 -0.07fF
C9 nCLK DFlipFlop_0/latch_diff_1/m1_657_280# 0.28fF
C10 nCLK DFlipFlop_1/latch_diff_1/nD 0.18fF
C11 nCLK DFlipFlop_2/latch_diff_1/nD 0.12fF
C12 sky130_fd_sc_hs__or2_1_0/a_152_368# Q1 0.01fF
C13 DFlipFlop_1/latch_diff_0/m1_657_280# CLK 0.31fF
C14 DFlipFlop_2/latch_diff_1/m1_657_280# Q2_d 0.03fF
C15 nCLK Q1 -0.02fF
C16 nCLK sky130_fd_sc_hs__or2_1_0/a_63_368# 0.05fF
C17 DFlipFlop_1/latch_diff_1/D CLK 0.18fF
C18 DFlipFlop_2/latch_diff_1/D Q2 0.13fF
C19 sky130_fd_sc_hs__or2_1_0/X nCLK_23 0.07fF
C20 DFlipFlop_1/D sky130_fd_sc_hs__or2_1_0/X 0.35fF
C21 DFlipFlop_2/latch_diff_1/D Q2_d 0.03fF
C22 sky130_fd_sc_hs__or2_1_1/X MC 0.02fF
C23 nCLK DFlipFlop_1/latch_diff_1/D 0.09fF
C24 vdd Q1 0.07fF
C25 Q2 DFlipFlop_2/nQ 0.13fF
C26 nCLK_23 sky130_fd_sc_hs__mux2_1_0/a_443_74# 0.09fF
C27 sky130_fd_sc_hs__or2_1_1/a_63_368# Q2 0.09fF
C28 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in CLK -0.10fF
C29 nCLK_23 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.49fF
C30 MC CLK 0.08fF
C31 nCLK_23 Q1 0.02fF
C32 DFlipFlop_0/nQ CLK 0.15fF
C33 DFlipFlop_2/latch_diff_1/nD Q2 0.17fF
C34 nCLK DFlipFlop_2/latch_diff_0/nD 0.09fF
C35 sky130_fd_sc_hs__or2_1_1/X vdd 0.03fF
C36 nCLK MC 0.01fF
C37 DFlipFlop_0/nQ nCLK 0.11fF
C38 vdd DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in 0.03fF
C39 sky130_fd_sc_hs__and2_1_0/a_56_136# CLK 0.08fF
C40 nCLK sky130_fd_sc_hs__or2_1_0/a_152_368# 0.01fF
C41 nCLK_23 sky130_fd_sc_hs__or2_1_1/X 0.26fF
C42 MC vdd 0.88fF
C43 vdd CLK 0.34fF
C44 CLK DFlipFlop_2/latch_diff_0/D 0.13fF
C45 sky130_fd_sc_hs__or2_1_1/X Q2 0.24fF
C46 sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__mux2_1_0/a_304_74# 0.08fF
C47 sky130_fd_sc_hs__or2_1_1/X Q2_d 0.03fF
C48 nCLK_23 MC 4.46fF
C49 nCLK vdd -0.55fF
C50 nCLK_23 DFlipFlop_0/nQ 0.05fF
C51 Q2 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in 0.38fF
C52 nCLK_23 CLK 0.22fF
C53 DFlipFlop_1/D CLK 0.40fF
C54 MC sky130_fd_sc_hs__mux2_1_0/a_27_112# 0.24fF
C55 MC Q2 0.18fF
C56 sky130_fd_sc_hs__mux2_1_0/a_524_368# nCLK_23 0.04fF
C57 DFlipFlop_0/latch_diff_1/nD Q1 0.03fF
C58 Q2 CLK 0.29fF
C59 CLK DFlipFlop_0/latch_diff_1/D 0.04fF
C60 nCLK_23 nCLK 0.11fF
C61 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out CLK 0.16fF
C62 DFlipFlop_0/latch_diff_0/m1_657_280# CLK 0.29fF
C63 DFlipFlop_0/latch_diff_0/nD nCLK_23 0.12fF
C64 DFlipFlop_1/D nCLK 0.16fF
C65 nCLK DFlipFlop_1/latch_diff_1/m1_657_280# 0.31fF
C66 nCLK_23 sky130_fd_sc_hs__and2_1_0/a_56_136# 0.14fF
C67 nCLK Q2 0.29fF
C68 sky130_fd_sc_hs__or2_1_0/X Q1 0.06fF
C69 nCLK_23 vdd 3.35fF
C70 vdd CLK_23 0.16fF
C71 DFlipFlop_1/latch_diff_0/nD CLK 0.09fF
C72 DFlipFlop_2/latch_diff_0/m1_657_280# nCLK 0.31fF
C73 nCLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in -0.02fF
C74 DFlipFlop_1/D vdd 0.07fF
C75 vdd Q2 1.63fF
C76 Q2 DFlipFlop_2/latch_diff_0/D 0.30fF
C77 DFlipFlop_0/latch_diff_1/m1_657_280# Q1 0.06fF
C78 vdd Q2_d 0.02fF
C79 sky130_fd_sc_hs__and2_1_0/a_143_136# nCLK_23 0.02fF
C80 nCLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out 0.06fF
C81 DFlipFlop_1/D nCLK_23 0.02fF
C82 nCLK_23 sky130_fd_sc_hs__mux2_1_0/a_27_112# 0.07fF
C83 nCLK_23 Q2 0.03fF
C84 DFlipFlop_0/latch_diff_1/nD CLK 0.02fF
C85 nCLK_23 DFlipFlop_0/latch_diff_1/D 0.05fF
C86 DFlipFlop_2/latch_diff_1/m1_657_280# CLK 0.33fF
C87 sky130_fd_sc_hs__or2_1_0/a_63_368# Q1 0.09fF
C88 nCLK_23 sky130_fd_sc_hs__mux2_1_0/a_304_74# 0.04fF
C89 CLK_23 sky130_fd_sc_hs__mux2_1_0/a_304_74# 0.05fF
C90 nCLK DFlipFlop_1/latch_diff_0/D 0.02fF
C91 vdd DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C92 DFlipFlop_2/latch_diff_1/D CLK 0.09fF
C93 nCLK DFlipFlop_0/latch_diff_1/nD 0.05fF
C94 sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__mux2_1_0/a_443_74# 0.03fF
C95 Q2 Q2_d 0.66fF
C96 sky130_fd_sc_hs__or2_1_0/X MC 0.09fF
C97 sky130_fd_sc_hs__or2_1_0/X CLK 0.01fF
C98 nCLK DFlipFlop_2/latch_diff_1/D 0.16fF
C99 DFlipFlop_2/nQ CLK 0.02fF
C100 sky130_fd_sc_hs__or2_1_0/X nCLK 0.06fF
C101 sky130_fd_sc_hs__or2_1_1/a_63_368# vss 0.37fF
C102 sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C103 sky130_fd_sc_hs__or2_1_0/X vss 0.92fF
C104 sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.39fF
C105 DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.72fF
C106 DFlipFlop_1/latch_diff_1/D vss -1.72fF
C107 DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C108 DFlipFlop_1/latch_diff_1/nD vss 0.58fF
C109 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C110 DFlipFlop_1/latch_diff_0/D vss 0.96fF
C111 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C112 DFlipFlop_1/D vss 2.98fF
C113 DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C114 Q2_d vss -0.22fF
C115 DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C116 DFlipFlop_2/nQ vss 0.48fF
C117 DFlipFlop_2/latch_diff_1/D vss -1.73fF
C118 DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C119 DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C120 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.94fF
C121 DFlipFlop_2/latch_diff_0/D vss 0.96fF
C122 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.84fF
C123 Q2 vss 1.35fF
C124 DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C125 Q1 vss 0.50fF
C126 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C127 nCLK vss -1.49fF
C128 DFlipFlop_0/nQ vss 0.48fF
C129 DFlipFlop_0/latch_diff_1/D vss -1.73fF
C130 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C131 CLK vss -0.61fF
C132 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C133 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C134 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C135 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C136 nCLK_23 vss -0.65fF
C137 vdd vss 115.92fF
C138 DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C139 CLK_23 vss -0.57fF
C140 sky130_fd_sc_hs__or2_1_1/X vss -0.35fF
C141 MC vss 2.09fF
C142 sky130_fd_sc_hs__mux2_1_0/a_304_74# vss 0.41fF
C143 sky130_fd_sc_hs__mux2_1_0/a_27_112# vss 0.69fF
.ends

.subckt freq_div clk_0 vss in_a n_clk_0 vdd prescaler_23_0/Q2 s_0 s_1_n s_1 prescaler_23_0/nCLK_23
+ prescaler_23_0/MC clk_d prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# s_0_n
+ clk_pre div_by_5_0/DFlipFlop_2/latch_diff_0/nD prescaler_23_0/DFlipFlop_2/latch_diff_1/D
+ prescaler_23_0/DFlipFlop_2/latch_diff_1/nD clk_1 div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280#
+ clk_out_mux21 n_clk_1 out div_by_5_0/Q1 div_by_5_0/DFlipFlop_2/latch_diff_0/D prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280#
+ div_by_5_0/DFlipFlop_2/latch_diff_1/nD clk_2 in_b clk_5 prescaler_23_0/DFlipFlop_2/latch_diff_0/nD
+ div_by_5_0/DFlipFlop_2/latch_diff_1/D prescaler_23_0/DFlipFlop_2/latch_diff_0/D
Xdiv_by_2_0 vss vdd div_by_2_0/nout_div div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in
+ clk_2 div_by_2_0/nCLK_2 div_by_2_0/o1 clk_out_mux21 div_by_2_0/out_div div_by_2_0/o2
+ div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out div_by_2
Xmux2to1_0 vss s_0_n clk_out_mux21 clk_pre clk_5 s_0 vdd mux2to1
Xinverter_min_x4_0 vdd inverter_min_x4_0/in vss clk_d inverter_min_x4
Xmux2to1_1 vss s_1_n out clk_d clk_2 s_1 vdd mux2to1
Xinverter_min_x2_0 clk_out_mux21 inverter_min_x4_0/in vss vdd inverter_min_x2
Xinverter_min_x2_1 s_1 s_1_n vss vdd inverter_min_x2
Xinverter_min_x2_2 s_0 s_0_n vss vdd inverter_min_x2
Xdiv_by_5_0 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in n_clk_1 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in
+ div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss vdd div_by_5_0/DFlipFlop_2/latch_diff_0/nD
+ div_by_5_0/Q0 div_by_5_0/Q1 clk_1 div_by_5_0/DFlipFlop_0/Q div_by_5_0/DFlipFlop_2/latch_diff_1/D
+ div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136#
+ div_by_5_0/nQ0 div_by_5_0/DFlipFlop_3/latch_diff_0/D div_by_5_0/DFlipFlop_3/latch_diff_1/nD
+ div_by_5_0/DFlipFlop_1/latch_diff_1/nD div_by_5_0/DFlipFlop_1/latch_diff_0/nD div_by_5_0/DFlipFlop_1/latch_diff_0/D
+ div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# clk_5 div_by_5_0/Q1_shift div_by_5_0/nQ2
+ div_by_5_0/DFlipFlop_2/D div_by_5_0/DFlipFlop_2/latch_diff_1/nD div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_1/latch_diff_1/D div_by_5_0/DFlipFlop_1/D div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ div_by_5_0/DFlipFlop_0/latch_diff_0/nD div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368#
+ div_by_5_0/DFlipFlop_0/D div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_0/latch_diff_1/D div_by_5_0/DFlipFlop_2/nQ div_by_5_0/DFlipFlop_3/latch_diff_0/nD
+ div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out div_by_5_0/DFlipFlop_2/latch_diff_0/D
+ div_by_5_0/DFlipFlop_0/latch_diff_0/D div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ div_by_5_0/DFlipFlop_3/latch_diff_1/D div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368#
+ div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136#
+ div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_152_368# div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# div_by_5_0/DFlipFlop_3/nQ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136#
+ div_by_5
Xmux2to4_0 vss n_clk_1 vdd s_0 s_0_n in_a clk_0 clk_1 n_clk_0 in_b mux2to4
Xprescaler_23_0 n_clk_0 vss prescaler_23_0/DFlipFlop_0/latch_diff_1/nD prescaler_23_0/nCLK_23
+ prescaler_23_0/DFlipFlop_2/latch_diff_0/nD vdd prescaler_23_0/DFlipFlop_2/latch_diff_1/D
+ prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out clk_pre prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280#
+ clk_0 prescaler_23_0/DFlipFlop_2/latch_diff_1/nD prescaler_23_0/DFlipFlop_0/latch_diff_0/nD
+ prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# prescaler_23_0/DFlipFlop_0/latch_diff_1/D
+ prescaler_23_0/DFlipFlop_2/latch_diff_0/D prescaler_23_0/MC prescaler_23_0/DFlipFlop_0/latch_diff_0/D
+ prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in prescaler_23_0/Q2
+ prescaler_23
C0 clk_pre prescaler_23_0/nCLK_23 0.03fF
C1 div_by_5_0/DFlipFlop_2/latch_diff_1/D s_0 0.05fF
C2 vdd s_0 3.90fF
C3 in_a clk_1 0.05fF
C4 clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_1/nD 0.09fF
C5 s_0_n div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# 0.05fF
C6 s_0_n div_by_5_0/DFlipFlop_1/latch_diff_1/nD 0.24fF
C7 vdd clk_5 0.06fF
C8 s_0 div_by_5_0/DFlipFlop_1/latch_diff_1/D 0.05fF
C9 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out s_0 0.30fF
C10 s_0 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out -0.19fF
C11 in_b s_0_n 0.48fF
C12 s_0 div_by_5_0/nQ2 0.05fF
C13 in_a s_0 0.30fF
C14 clk_pre vdd 0.17fF
C15 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out s_0_n -0.01fF
C16 s_0_n clk_1 4.82fF
C17 div_by_5_0/DFlipFlop_0/D s_0_n 0.05fF
C18 vdd inverter_min_x4_0/in 0.09fF
C19 s_0_n s_0 7.76fF
C20 div_by_5_0/Q1 vdd 0.04fF
C21 n_clk_0 prescaler_23_0/nCLK_23 0.16fF
C22 s_0_n clk_5 0.56fF
C23 div_by_5_0/DFlipFlop_2/latch_diff_0/nD s_0_n 0.20fF
C24 div_by_5_0/DFlipFlop_2/nQ s_0 0.05fF
C25 n_clk_1 div_by_5_0/DFlipFlop_0/latch_diff_0/D 0.11fF
C26 n_clk_0 vdd 0.25fF
C27 clk_2 vdd 0.06fF
C28 s_1 clk_d 0.22fF
C29 clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_1/D 0.13fF
C30 div_by_5_0/Q1 s_0_n 0.21fF
C31 clk_out_mux21 s_0 0.68fF
C32 s_0 div_by_5_0/DFlipFlop_2/D 0.03fF
C33 div_by_5_0/DFlipFlop_3/latch_diff_0/D s_0 0.10fF
C34 vdd div_by_5_0/Q0 0.05fF
C35 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# n_clk_1 0.06fF
C36 clk_out_mux21 clk_5 0.05fF
C37 n_clk_1 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.11fF
C38 clk_pre clk_out_mux21 1.19fF
C39 n_clk_0 s_0_n 0.31fF
C40 div_by_5_0/DFlipFlop_2/latch_diff_1/nD s_0_n 0.24fF
C41 div_by_5_0/DFlipFlop_3/latch_diff_1/D s_0_n 0.24fF
C42 n_clk_1 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.14fF
C43 div_by_5_0/DFlipFlop_0/latch_diff_0/nD s_0_n 0.20fF
C44 div_by_5_0/Q1_shift s_0_n 0.04fF
C45 div_by_5_0/Q1_shift div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_152_368# -0.02fF
C46 in_b n_clk_1 0.05fF
C47 s_0_n div_by_5_0/Q0 0.24fF
C48 div_by_5_0/nQ0 s_0 0.05fF
C49 div_by_5_0/DFlipFlop_3/latch_diff_1/nD s_0 0.05fF
C50 div_by_5_0/DFlipFlop_0/D n_clk_1 0.21fF
C51 div_by_5_0/DFlipFlop_3/nQ s_0 0.02fF
C52 s_0 div_by_5_0/DFlipFlop_1/latch_diff_0/nD 0.12fF
C53 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in s_0 -0.36fF
C54 n_clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_1/nD 0.13fF
C55 s_0_n div_by_5_0/DFlipFlop_1/D 0.19fF
C56 s_0 div_by_5_0/DFlipFlop_0/Q 0.02fF
C57 s_1 out 0.39fF
C58 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# n_clk_1 0.03fF
C59 s_0_n div_by_5_0/DFlipFlop_0/latch_diff_1/D 0.04fF
C60 clk_d inverter_min_x4_0/in 0.11fF
C61 div_by_5_0/DFlipFlop_0/latch_diff_1/nD clk_1 0.08fF
C62 div_by_5_0/DFlipFlop_2/latch_diff_1/D s_0_n 0.04fF
C63 s_0_n vdd 2.76fF
C64 s_0 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.02fF
C65 s_1 s_1_n 0.39fF
C66 n_clk_1 div_by_5_0/Q1 0.15fF
C67 s_0_n div_by_5_0/DFlipFlop_1/latch_diff_1/D 0.04fF
C68 s_0_n div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out 0.31fF
C69 s_0_n div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out -0.29fF
C70 s_0_n div_by_5_0/nQ2 0.05fF
C71 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out clk_1 0.05fF
C72 s_0 div_by_5_0/DFlipFlop_1/latch_diff_1/nD 0.02fF
C73 div_by_5_0/DFlipFlop_0/D clk_1 0.14fF
C74 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out s_0 -0.13fF
C75 s_0 clk_1 1.36fF
C76 prescaler_23_0/DFlipFlop_0/latch_diff_1/D n_clk_0 0.09fF
C77 div_by_5_0/DFlipFlop_0/D s_0 0.03fF
C78 clk_out_mux21 vdd 0.14fF
C79 out s_1_n 0.33fF
C80 div_by_5_0/DFlipFlop_2/nQ s_0_n 0.04fF
C81 n_clk_1 div_by_5_0/Q0 0.01fF
C82 div_by_5_0/Q1 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in -0.03fF
C83 div_by_5_0/DFlipFlop_2/latch_diff_0/nD s_0 0.12fF
C84 clk_pre s_0 0.21fF
C85 clk_0 prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.16fF
C86 clk_out_mux21 s_0_n 0.45fF
C87 s_0_n div_by_5_0/DFlipFlop_2/D 0.05fF
C88 s_0_n div_by_5_0/DFlipFlop_3/latch_diff_0/D 0.17fF
C89 n_clk_1 div_by_5_0/DFlipFlop_0/latch_diff_1/D 0.08fF
C90 div_by_5_0/Q1 s_0 0.04fF
C91 clk_0 prescaler_23_0/nCLK_23 0.16fF
C92 vdd clk_d 0.23fF
C93 n_clk_0 clk_1 -0.03fF
C94 n_clk_1 vdd 0.15fF
C95 clk_2 out 0.05fF
C96 clk_0 vdd 0.63fF
C97 div_by_5_0/DFlipFlop_2/latch_diff_1/nD s_0 0.02fF
C98 div_by_5_0/DFlipFlop_0/latch_diff_0/nD clk_1 0.08fF
C99 clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_0/nD 0.09fF
C100 div_by_5_0/DFlipFlop_3/latch_diff_1/D s_0 0.02fF
C101 div_by_5_0/nQ0 s_0_n 0.05fF
C102 div_by_5_0/DFlipFlop_0/latch_diff_0/nD s_0 0.12fF
C103 div_by_5_0/Q1_shift s_0 0.05fF
C104 clk_2 s_1_n 0.59fF
C105 div_by_5_0/DFlipFlop_3/latch_diff_1/nD s_0_n 0.04fF
C106 s_0_n div_by_5_0/DFlipFlop_3/nQ 0.24fF
C107 s_0 div_by_5_0/Q0 0.02fF
C108 div_by_5_0/Q1_shift clk_5 0.04fF
C109 s_0_n div_by_5_0/DFlipFlop_1/latch_diff_0/nD 0.20fF
C110 s_0_n div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in -0.37fF
C111 n_clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_0/D 0.13fF
C112 s_0_n div_by_5_0/DFlipFlop_0/Q 0.24fF
C113 clk_1 div_by_5_0/DFlipFlop_0/latch_diff_1/D 0.11fF
C114 s_0 div_by_5_0/DFlipFlop_1/D 0.03fF
C115 n_clk_0 prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.14fF
C116 s_0 div_by_5_0/DFlipFlop_0/latch_diff_1/D 0.05fF
C117 vdd clk_1 0.18fF
C118 s_0_n div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.24fF
C119 prescaler_23_0/sky130_fd_sc_hs__or2_1_1/a_63_368# vss 0.37fF
C120 prescaler_23_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C121 prescaler_23_0/sky130_fd_sc_hs__or2_1_0/X vss 0.49fF
C122 prescaler_23_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C123 prescaler_23_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C124 prescaler_23_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C125 prescaler_23_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C126 prescaler_23_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C127 prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C128 prescaler_23_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C129 prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C130 prescaler_23_0/DFlipFlop_1/D vss 1.90fF
C131 prescaler_23_0/DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C132 prescaler_23_0/Q2_d vss -0.69fF
C133 prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C134 prescaler_23_0/DFlipFlop_2/nQ vss 0.48fF
C135 prescaler_23_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C136 prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C137 prescaler_23_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C138 prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C139 prescaler_23_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C140 prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C141 prescaler_23_0/Q2 vss 0.55fF
C142 prescaler_23_0/DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C143 prescaler_23_0/Q1 vss 0.07fF
C144 prescaler_23_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C145 n_clk_0 vss -5.72fF
C146 prescaler_23_0/DFlipFlop_0/nQ vss 0.48fF
C147 prescaler_23_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C148 prescaler_23_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C149 clk_0 vss 0.74fF
C150 prescaler_23_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C151 prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C152 prescaler_23_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C153 prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C154 prescaler_23_0/nCLK_23 vss -1.02fF
C155 prescaler_23_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C156 prescaler_23_0/sky130_fd_sc_hs__or2_1_1/X vss -1.01fF
C157 prescaler_23_0/MC vss 1.07fF
C158 prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_304_74# vss 0.36fF
C159 prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_27_112# vss 0.65fF
C160 in_b vss 2.26fF
C161 s_0_n vss -2.65fF
C162 in_a vss 2.25fF
C163 s_0 vss 5.73fF
C164 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C165 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.38fF
C166 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C167 div_by_5_0/Q1_shift vss -0.36fF
C168 div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.57fF
C169 div_by_5_0/DFlipFlop_3/nQ vss 0.48fF
C170 div_by_5_0/DFlipFlop_3/latch_diff_1/D vss -1.73fF
C171 div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C172 div_by_5_0/DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C173 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C174 div_by_5_0/DFlipFlop_3/latch_diff_0/D vss 0.96fF
C175 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C176 div_by_5_0/DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C177 div_by_5_0/Q1 vss 4.35fF
C178 div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C179 div_by_5_0/DFlipFlop_2/nQ vss 0.48fF
C180 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C181 div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C182 div_by_5_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C183 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C184 div_by_5_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C185 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C186 div_by_5_0/DFlipFlop_2/D vss 3.13fF
C187 div_by_5_0/DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C188 div_by_5_0/Q0 vss 0.29fF
C189 div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C190 div_by_5_0/nQ0 vss 0.99fF
C191 div_by_5_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C192 div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C193 div_by_5_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C194 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C195 div_by_5_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C196 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C197 div_by_5_0/DFlipFlop_1/D vss 3.64fF
C198 div_by_5_0/DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C199 div_by_5_0/DFlipFlop_0/Q vss -0.94fF
C200 div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C201 n_clk_1 vss -0.44fF
C202 div_by_5_0/nQ2 vss 1.38fF
C203 div_by_5_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C204 div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C205 clk_1 vss -1.17fF
C206 div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C207 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C208 div_by_5_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C209 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C210 div_by_5_0/DFlipFlop_0/D vss 3.96fF
C211 vdd vss 355.84fF
C212 div_by_5_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C213 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C214 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.40fF
C215 s_1_n vss 1.15fF
C216 out vss 1.17fF
C217 clk_d vss 0.79fF
C218 s_1 vss 2.97fF
C219 inverter_min_x4_0/in vss 2.77fF
C220 clk_5 vss 0.10fF
C221 clk_out_mux21 vss 5.62fF
C222 clk_pre vss 1.31fF
C223 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C224 div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C225 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C226 div_by_2_0/DFlipFlop_0/nCLK vss 1.03fF
C227 clk_2 vss 3.57fF
C228 div_by_2_0/o1 vss 2.20fF
C229 div_by_2_0/nCLK_2 vss 1.04fF
C230 div_by_2_0/o2 vss 2.08fF
C231 div_by_2_0/out_div vss -0.80fF
C232 div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C233 div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C234 div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C235 div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C236 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C237 div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C238 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C239 div_by_2_0/nout_div vss 2.62fF
C240 div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
.ends

.subckt sky130_fd_pr__nfet_01v8_CBAU6Y a_n73_n150# a_n33_n238# w_n211_n360# a_15_n150#
X0 a_15_n150# a_n33_n238# a_n73_n150# w_n211_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_15_n150# a_n33_n238# 0.02fF
C1 a_n73_n150# a_n33_n238# 0.02fF
C2 a_15_n150# a_n73_n150# 0.51fF
C3 a_15_n150# w_n211_n360# 0.23fF
C4 a_n73_n150# w_n211_n360# 0.23fF
C5 a_n33_n238# w_n211_n360# 0.17fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4757AC VSUBS a_n73_n150# a_n33_181# w_n211_n369# a_15_n150#
X0 a_15_n150# a_n33_181# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_15_n150# w_n211_n369# 0.20fF
C1 a_n73_n150# a_15_n150# 0.51fF
C2 a_n33_181# a_15_n150# 0.01fF
C3 a_n73_n150# w_n211_n369# 0.20fF
C4 a_n33_181# w_n211_n369# 0.05fF
C5 a_n73_n150# a_n33_181# 0.01fF
C6 a_15_n150# VSUBS 0.03fF
C7 a_n73_n150# VSUBS 0.03fF
C8 a_n33_181# VSUBS 0.13fF
C9 w_n211_n369# VSUBS 1.98fF
.ends

.subckt sky130_fd_pr__nfet_01v8_7H8F5S a_n465_172# a_n417_n150# a_351_n150# a_255_n150#
+ w_n647_n360# a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150#
X0 a_159_n150# a_n465_172# a_63_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n225_n150# a_n465_172# a_n321_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_447_n150# a_n465_172# a_351_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_63_n150# a_n465_172# a_n33_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n465_172# a_n225_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n465_172# a_n509_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n33_n150# a_n465_172# a_n129_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_351_n150# a_n465_172# a_255_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_255_n150# a_n465_172# a_159_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n321_n150# a_n465_172# a_n417_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_351_n150# a_255_n150# 0.43fF
C1 a_n129_n150# a_n465_172# 0.10fF
C2 a_n321_n150# a_63_n150# 0.07fF
C3 a_n321_n150# a_n465_172# 0.10fF
C4 a_n33_n150# a_n417_n150# 0.07fF
C5 a_447_n150# a_159_n150# 0.10fF
C6 a_447_n150# a_255_n150# 0.16fF
C7 a_n129_n150# a_n417_n150# 0.10fF
C8 a_n129_n150# a_n509_n150# 0.07fF
C9 a_n33_n150# a_n225_n150# 0.16fF
C10 a_n465_172# a_63_n150# 0.10fF
C11 a_n129_n150# a_n225_n150# 0.43fF
C12 a_n417_n150# a_n321_n150# 0.43fF
C13 a_n509_n150# a_n321_n150# 0.16fF
C14 a_447_n150# a_351_n150# 0.43fF
C15 a_n321_n150# a_n225_n150# 0.43fF
C16 a_n33_n150# a_159_n150# 0.16fF
C17 a_n33_n150# a_255_n150# 0.10fF
C18 a_n129_n150# a_159_n150# 0.10fF
C19 a_n129_n150# a_255_n150# 0.07fF
C20 a_n225_n150# a_63_n150# 0.10fF
C21 a_n417_n150# a_n465_172# 0.10fF
C22 a_n509_n150# a_n465_172# 0.01fF
C23 a_n33_n150# a_351_n150# 0.07fF
C24 a_n465_172# a_n225_n150# 0.10fF
C25 a_63_n150# a_159_n150# 0.43fF
C26 a_255_n150# a_63_n150# 0.16fF
C27 a_n417_n150# a_n509_n150# 0.43fF
C28 a_n465_172# a_159_n150# 0.10fF
C29 a_n465_172# a_255_n150# 0.10fF
C30 a_n417_n150# a_n225_n150# 0.16fF
C31 a_n509_n150# a_n225_n150# 0.10fF
C32 a_351_n150# a_63_n150# 0.10fF
C33 a_351_n150# a_n465_172# 0.10fF
C34 a_n33_n150# a_n129_n150# 0.43fF
C35 a_n225_n150# a_159_n150# 0.07fF
C36 a_447_n150# a_63_n150# 0.07fF
C37 a_n33_n150# a_n321_n150# 0.10fF
C38 a_447_n150# a_n465_172# 0.01fF
C39 a_n129_n150# a_n321_n150# 0.16fF
C40 a_255_n150# a_159_n150# 0.43fF
C41 a_n33_n150# a_63_n150# 0.43fF
C42 a_n129_n150# a_63_n150# 0.16fF
C43 a_n33_n150# a_n465_172# 0.10fF
C44 a_351_n150# a_159_n150# 0.16fF
C45 a_447_n150# w_n647_n360# 0.17fF
C46 a_351_n150# w_n647_n360# 0.10fF
C47 a_255_n150# w_n647_n360# 0.08fF
C48 a_159_n150# w_n647_n360# 0.07fF
C49 a_63_n150# w_n647_n360# 0.04fF
C50 a_n33_n150# w_n647_n360# 0.04fF
C51 a_n129_n150# w_n647_n360# 0.04fF
C52 a_n225_n150# w_n647_n360# 0.07fF
C53 a_n321_n150# w_n647_n360# 0.08fF
C54 a_n417_n150# w_n647_n360# 0.10fF
C55 a_n509_n150# w_n647_n360# 0.17fF
C56 a_n465_172# w_n647_n360# 1.49fF
.ends

.subckt sky130_fd_pr__pfet_01v8_8DL6ZL VSUBS a_n417_n150# a_351_n150# a_255_n150#
+ a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n465_n247# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150# w_n647_n369#
X0 a_63_n150# a_n465_n247# a_n33_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n129_n150# a_n465_n247# a_n225_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n417_n150# a_n465_n247# a_n509_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n33_n150# a_n465_n247# a_n129_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_351_n150# a_n465_n247# a_255_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_255_n150# a_n465_n247# a_159_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n321_n150# a_n465_n247# a_n417_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_159_n150# a_n465_n247# a_63_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n225_n150# a_n465_n247# a_n321_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_447_n150# a_n465_n247# a_351_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_63_n150# a_255_n150# 0.16fF
C1 a_159_n150# w_n647_n369# 0.04fF
C2 a_n465_n247# a_159_n150# 0.08fF
C3 a_n129_n150# a_n33_n150# 0.43fF
C4 a_n129_n150# a_63_n150# 0.16fF
C5 a_n225_n150# a_n33_n150# 0.16fF
C6 a_n417_n150# w_n647_n369# 0.07fF
C7 a_n417_n150# a_n465_n247# 0.08fF
C8 a_n225_n150# a_63_n150# 0.10fF
C9 a_255_n150# w_n647_n369# 0.05fF
C10 a_n465_n247# a_255_n150# 0.08fF
C11 a_n129_n150# w_n647_n369# 0.02fF
C12 a_n129_n150# a_n465_n247# 0.08fF
C13 a_n417_n150# a_n509_n150# 0.43fF
C14 a_n225_n150# w_n647_n369# 0.04fF
C15 a_n225_n150# a_n465_n247# 0.08fF
C16 a_159_n150# a_255_n150# 0.43fF
C17 a_n321_n150# a_n33_n150# 0.10fF
C18 a_n509_n150# a_n129_n150# 0.07fF
C19 a_n321_n150# a_63_n150# 0.07fF
C20 a_n129_n150# a_159_n150# 0.10fF
C21 a_351_n150# a_447_n150# 0.43fF
C22 a_351_n150# a_n33_n150# 0.07fF
C23 a_n509_n150# a_n225_n150# 0.10fF
C24 a_351_n150# a_63_n150# 0.10fF
C25 a_n225_n150# a_159_n150# 0.07fF
C26 a_n417_n150# a_n129_n150# 0.10fF
C27 a_63_n150# a_447_n150# 0.07fF
C28 a_63_n150# a_n33_n150# 0.43fF
C29 a_n417_n150# a_n225_n150# 0.16fF
C30 a_n129_n150# a_255_n150# 0.07fF
C31 a_n321_n150# w_n647_n369# 0.05fF
C32 a_n321_n150# a_n465_n247# 0.08fF
C33 a_351_n150# w_n647_n369# 0.07fF
C34 a_351_n150# a_n465_n247# 0.08fF
C35 a_447_n150# w_n647_n369# 0.14fF
C36 a_n33_n150# w_n647_n369# 0.02fF
C37 a_n225_n150# a_n129_n150# 0.43fF
C38 a_n465_n247# a_n33_n150# 0.08fF
C39 a_n509_n150# a_n321_n150# 0.16fF
C40 a_63_n150# w_n647_n369# 0.02fF
C41 a_63_n150# a_n465_n247# 0.08fF
C42 a_351_n150# a_159_n150# 0.16fF
C43 a_n417_n150# a_n321_n150# 0.43fF
C44 a_447_n150# a_159_n150# 0.10fF
C45 a_n33_n150# a_159_n150# 0.16fF
C46 a_n465_n247# w_n647_n369# 0.47fF
C47 a_63_n150# a_159_n150# 0.43fF
C48 a_n417_n150# a_n33_n150# 0.07fF
C49 a_351_n150# a_255_n150# 0.43fF
C50 a_n129_n150# a_n321_n150# 0.16fF
C51 a_447_n150# a_255_n150# 0.16fF
C52 a_n33_n150# a_255_n150# 0.10fF
C53 a_n225_n150# a_n321_n150# 0.43fF
C54 a_n509_n150# w_n647_n369# 0.14fF
C55 a_447_n150# VSUBS 0.03fF
C56 a_351_n150# VSUBS 0.03fF
C57 a_255_n150# VSUBS 0.03fF
C58 a_159_n150# VSUBS 0.03fF
C59 a_63_n150# VSUBS 0.03fF
C60 a_n33_n150# VSUBS 0.03fF
C61 a_n129_n150# VSUBS 0.03fF
C62 a_n225_n150# VSUBS 0.03fF
C63 a_n321_n150# VSUBS 0.03fF
C64 a_n417_n150# VSUBS 0.03fF
C65 a_n509_n150# VSUBS 0.03fF
C66 a_n465_n247# VSUBS 1.07fF
C67 w_n647_n369# VSUBS 4.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EDT3AT a_15_n11# a_n33_n99# w_n211_n221# a_n73_n11#
X0 a_15_n11# a_n33_n99# a_n73_n11# w_n211_n221# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n33_n99# a_15_n11# 0.02fF
C1 a_n73_n11# a_15_n11# 0.15fF
C2 a_n33_n99# a_n73_n11# 0.02fF
C3 a_15_n11# w_n211_n221# 0.09fF
C4 a_n73_n11# w_n211_n221# 0.09fF
C5 a_n33_n99# w_n211_n221# 0.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AQR2CW a_n33_66# a_n78_n106# w_n216_n254# a_20_n106#
X0 a_20_n106# a_n33_66# a_n78_n106# w_n216_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=200000u
C0 a_n78_n106# a_20_n106# 0.21fF
C1 a_20_n106# w_n216_n254# 0.14fF
C2 a_n78_n106# w_n216_n254# 0.14fF
C3 a_n33_66# w_n216_n254# 0.12fF
.ends

.subckt sky130_fd_pr__pfet_01v8_HRYSXS VSUBS a_n33_n211# a_n78_n114# w_n216_n334#
+ a_20_n114#
X0 a_20_n114# a_n33_n211# a_n78_n114# w_n216_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=200000u
C0 w_n216_n334# a_n78_n114# 0.20fF
C1 a_20_n114# w_n216_n334# 0.20fF
C2 a_20_n114# a_n78_n114# 0.42fF
C3 a_20_n114# VSUBS 0.03fF
C4 a_n78_n114# VSUBS 0.03fF
C5 a_n33_n211# VSUBS 0.12fF
C6 w_n216_n334# VSUBS 1.66fF
.ends

.subckt inverter_csvco in vbulkn out vbulkp vdd vss
Xsky130_fd_pr__nfet_01v8_AQR2CW_0 in vss vbulkn out sky130_fd_pr__nfet_01v8_AQR2CW
Xsky130_fd_pr__pfet_01v8_HRYSXS_0 vbulkn in vdd vbulkp out sky130_fd_pr__pfet_01v8_HRYSXS
C0 in vss 0.01fF
C1 vbulkp vdd 0.04fF
C2 vbulkp out 0.08fF
C3 in vdd 0.01fF
C4 in out 0.11fF
C5 vbulkp vbulkn 2.49fF
C6 out vbulkn 0.60fF
C7 vdd vbulkn 0.06fF
C8 in vbulkn 0.54fF
C9 vss vbulkn 0.17fF
.ends

.subckt csvco_branch vctrl inverter_csvco_0/vdd in vbp cap_vco_0/t D0 vss out vdd
+ inverter_csvco_0/vss
Xsky130_fd_pr__nfet_01v8_7H8F5S_0 vctrl inverter_csvco_0/vss inverter_csvco_0/vss
+ vss vss inverter_csvco_0/vss vss vss inverter_csvco_0/vss vss inverter_csvco_0/vss
+ vss vss sky130_fd_pr__nfet_01v8_7H8F5S
Xsky130_fd_pr__pfet_01v8_8DL6ZL_0 vss inverter_csvco_0/vdd inverter_csvco_0/vdd vdd
+ inverter_csvco_0/vdd vdd vdd inverter_csvco_0/vdd vbp vdd inverter_csvco_0/vdd vdd
+ vdd vdd sky130_fd_pr__pfet_01v8_8DL6ZL
Xsky130_fd_pr__nfet_01v8_EDT3AT_0 cap_vco_0/t D0 vss out sky130_fd_pr__nfet_01v8_EDT3AT
Xinverter_csvco_0 in vss out vdd inverter_csvco_0/vdd inverter_csvco_0/vss inverter_csvco
C0 inverter_csvco_0/vdd cap_vco_0/t 0.10fF
C1 D0 out 0.09fF
C2 vdd cap_vco_0/t 0.04fF
C3 in out 0.06fF
C4 out inverter_csvco_0/vdd 0.02fF
C5 out inverter_csvco_0/vss 0.03fF
C6 vbp inverter_csvco_0/vdd 0.75fF
C7 in inverter_csvco_0/vdd 0.01fF
C8 vbp vdd 1.21fF
C9 D0 inverter_csvco_0/vss 0.02fF
C10 vctrl inverter_csvco_0/vss 0.87fF
C11 inverter_csvco_0/vdd vdd 1.89fF
C12 in inverter_csvco_0/vss 0.01fF
C13 out cap_vco_0/t 0.70fF
C14 out vss 0.93fF
C15 inverter_csvco_0/vdd vss 0.26fF
C16 in vss 0.69fF
C17 D0 vss -0.67fF
C18 vbp vss 0.13fF
C19 vdd vss 9.58fF
C20 cap_vco_0/t vss 7.22fF
C21 inverter_csvco_0/vss vss 1.79fF
C22 vctrl vss 3.06fF
.ends

.subckt ring_osc csvco_branch_0/inverter_csvco_0/vdd vctrl vss csvco_branch_1/inverter_csvco_0/vdd
+ csvco_branch_2/inverter_csvco_0/vdd vdd csvco_branch_2/vbp csvco_branch_0/inverter_csvco_0/vss
+ D0 csvco_branch_2/cap_vco_0/t out_vco
Xsky130_fd_pr__nfet_01v8_CBAU6Y_0 vss vctrl vss csvco_branch_2/vbp sky130_fd_pr__nfet_01v8_CBAU6Y
Xsky130_fd_pr__pfet_01v8_4757AC_0 vss vdd csvco_branch_2/vbp vdd csvco_branch_2/vbp
+ sky130_fd_pr__pfet_01v8_4757AC
Xcsvco_branch_0 vctrl csvco_branch_0/inverter_csvco_0/vdd out_vco csvco_branch_2/vbp
+ csvco_branch_0/cap_vco_0/t D0 vss csvco_branch_1/in vdd csvco_branch_0/inverter_csvco_0/vss
+ csvco_branch
Xcsvco_branch_2 vctrl csvco_branch_2/inverter_csvco_0/vdd csvco_branch_2/in csvco_branch_2/vbp
+ csvco_branch_2/cap_vco_0/t D0 vss out_vco vdd csvco_branch_2/inverter_csvco_0/vss
+ csvco_branch
Xcsvco_branch_1 vctrl csvco_branch_1/inverter_csvco_0/vdd csvco_branch_1/in csvco_branch_2/vbp
+ csvco_branch_1/cap_vco_0/t D0 vss csvco_branch_2/in vdd csvco_branch_1/inverter_csvco_0/vss
+ csvco_branch
C0 csvco_branch_0/inverter_csvco_0/vdd csvco_branch_2/vbp 0.06fF
C1 vctrl csvco_branch_2/vbp 0.06fF
C2 out_vco csvco_branch_0/cap_vco_0/t 0.03fF
C3 csvco_branch_0/inverter_csvco_0/vss csvco_branch_2/vbp 0.06fF
C4 csvco_branch_1/inverter_csvco_0/vss D0 0.68fF
C5 vdd csvco_branch_1/inverter_csvco_0/vdd 0.19fF
C6 out_vco csvco_branch_2/in 0.58fF
C7 csvco_branch_0/inverter_csvco_0/vdd vdd 0.13fF
C8 csvco_branch_2/inverter_csvco_0/vss D0 0.68fF
C9 vdd csvco_branch_2/vbp 1.49fF
C10 csvco_branch_1/in out_vco 0.76fF
C11 out_vco csvco_branch_1/cap_vco_0/t 0.03fF
C12 D0 vctrl 4.41fF
C13 csvco_branch_2/inverter_csvco_0/vdd vdd 0.10fF
C14 csvco_branch_0/inverter_csvco_0/vss D0 0.49fF
C15 csvco_branch_2/in vss 1.60fF
C16 csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C17 csvco_branch_1/cap_vco_0/t vss 7.10fF
C18 csvco_branch_1/inverter_csvco_0/vss vss 0.72fF
C19 csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C20 csvco_branch_2/cap_vco_0/t vss 7.10fF
C21 csvco_branch_2/inverter_csvco_0/vss vss 0.62fF
C22 csvco_branch_1/in vss 1.58fF
C23 csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C24 out_vco vss 0.67fF
C25 D0 vss -1.55fF
C26 vdd vss 31.40fF
C27 csvco_branch_0/cap_vco_0/t vss 7.10fF
C28 csvco_branch_0/inverter_csvco_0/vss vss 0.66fF
C29 vctrl vss 11.02fF
C30 csvco_branch_2/vbp vss 0.77fF
.ends

.subckt ring_osc_buffer vss in_vco vdd o1 out_div out_pad
Xinverter_min_x4_1 vdd out_div vss out_pad inverter_min_x4
Xinverter_min_x4_0 vdd o1 vss out_div inverter_min_x4
Xinverter_min_x2_0 in_vco o1 vss vdd inverter_min_x2
C0 out_div o1 0.11fF
C1 out_div vdd 0.17fF
C2 vdd o1 0.09fF
C3 out_div out_pad 0.15fF
C4 vdd out_pad 0.10fF
C5 in_vco vss 0.83fF
C6 o1 vss 2.72fF
C7 vdd vss 14.54fF
C8 out_pad vss 0.70fF
C9 out_div vss 3.00fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AZESM8 a_n63_n151# a_n33_n125# a_n255_n151# a_33_n151#
+ a_n225_n125# a_63_n125# a_n129_n125# a_n159_n151# w_n455_n335# a_225_n151# a_255_n125#
+ a_129_n151# a_159_n125# a_n317_n125#
X0 a_159_n125# a_129_n151# a_63_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n225_n125# a_n255_n151# a_n317_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_63_n125# a_33_n151# a_n33_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_n129_n125# a_n159_n151# a_n225_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n33_n125# a_n63_n151# a_n129_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_255_n125# a_225_n151# a_159_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_33_n151# a_n63_n151# 0.02fF
C1 a_159_n125# a_n33_n125# 0.13fF
C2 a_129_n151# a_33_n151# 0.02fF
C3 a_n33_n125# a_n317_n125# 0.08fF
C4 a_159_n125# a_n129_n125# 0.08fF
C5 a_n159_n151# a_n63_n151# 0.02fF
C6 a_159_n125# a_63_n125# 0.36fF
C7 a_n317_n125# a_n129_n125# 0.13fF
C8 a_n317_n125# a_63_n125# 0.06fF
C9 a_159_n125# a_n225_n125# 0.06fF
C10 a_n317_n125# a_n225_n125# 0.36fF
C11 a_159_n125# a_255_n125# 0.36fF
C12 a_n33_n125# a_n129_n125# 0.36fF
C13 a_n33_n125# a_63_n125# 0.36fF
C14 a_n33_n125# a_n225_n125# 0.13fF
C15 a_n129_n125# a_63_n125# 0.13fF
C16 a_n129_n125# a_n225_n125# 0.36fF
C17 a_n225_n125# a_63_n125# 0.08fF
C18 a_255_n125# a_n33_n125# 0.08fF
C19 a_129_n151# a_225_n151# 0.02fF
C20 a_255_n125# a_n129_n125# 0.06fF
C21 a_255_n125# a_63_n125# 0.13fF
C22 a_n255_n151# a_n159_n151# 0.02fF
C23 a_255_n125# w_n455_n335# 0.14fF
C24 a_159_n125# w_n455_n335# 0.08fF
C25 a_63_n125# w_n455_n335# 0.07fF
C26 a_n33_n125# w_n455_n335# 0.08fF
C27 a_n129_n125# w_n455_n335# 0.07fF
C28 a_n225_n125# w_n455_n335# 0.08fF
C29 a_n317_n125# w_n455_n335# 0.14fF
C30 a_225_n151# w_n455_n335# 0.05fF
C31 a_129_n151# w_n455_n335# 0.05fF
C32 a_33_n151# w_n455_n335# 0.05fF
C33 a_n63_n151# w_n455_n335# 0.05fF
C34 a_n159_n151# w_n455_n335# 0.05fF
C35 a_n255_n151# w_n455_n335# 0.05fF
.ends

.subckt sky130_fd_pr__pfet_01v8_XJXT7S VSUBS a_n33_n125# a_n255_n154# a_33_n154# a_n225_n125#
+ a_n159_n154# a_63_n125# a_n129_n125# a_225_n154# a_129_n154# a_255_n125# a_159_n125#
+ a_n317_n125# w_n455_n344# a_n63_n154#
X0 a_n129_n125# a_n159_n154# a_n225_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n33_n125# a_n63_n154# a_n129_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_255_n125# a_225_n154# a_159_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_159_n125# a_129_n154# a_63_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n225_n125# a_n255_n154# a_n317_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_63_n125# a_33_n154# a_n33_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_159_n125# w_n455_n344# 0.06fF
C1 a_n225_n125# a_159_n125# 0.06fF
C2 w_n455_n344# a_63_n125# 0.04fF
C3 a_n225_n125# a_63_n125# 0.08fF
C4 a_n129_n125# w_n455_n344# 0.04fF
C5 a_n33_n125# w_n455_n344# 0.05fF
C6 a_n225_n125# a_n129_n125# 0.36fF
C7 a_n225_n125# a_n33_n125# 0.13fF
C8 a_255_n125# w_n455_n344# 0.11fF
C9 a_n317_n125# w_n455_n344# 0.11fF
C10 a_n225_n125# a_n317_n125# 0.36fF
C11 a_n63_n154# a_n159_n154# 0.02fF
C12 a_33_n154# a_129_n154# 0.02fF
C13 a_n63_n154# a_33_n154# 0.02fF
C14 a_159_n125# a_63_n125# 0.36fF
C15 a_n255_n154# a_n159_n154# 0.02fF
C16 a_159_n125# a_n129_n125# 0.08fF
C17 a_n33_n125# a_159_n125# 0.13fF
C18 a_255_n125# a_159_n125# 0.36fF
C19 a_n225_n125# w_n455_n344# 0.06fF
C20 a_n129_n125# a_63_n125# 0.13fF
C21 a_n33_n125# a_63_n125# 0.36fF
C22 a_255_n125# a_63_n125# 0.13fF
C23 a_n317_n125# a_63_n125# 0.06fF
C24 a_n33_n125# a_n129_n125# 0.36fF
C25 a_255_n125# a_n129_n125# 0.06fF
C26 a_255_n125# a_n33_n125# 0.08fF
C27 a_n129_n125# a_n317_n125# 0.13fF
C28 a_n33_n125# a_n317_n125# 0.08fF
C29 a_225_n154# a_129_n154# 0.02fF
C30 a_255_n125# VSUBS 0.03fF
C31 a_159_n125# VSUBS 0.03fF
C32 a_63_n125# VSUBS 0.03fF
C33 a_n33_n125# VSUBS 0.03fF
C34 a_n129_n125# VSUBS 0.03fF
C35 a_n225_n125# VSUBS 0.03fF
C36 a_n317_n125# VSUBS 0.03fF
C37 a_225_n154# VSUBS 0.05fF
C38 a_129_n154# VSUBS 0.05fF
C39 a_33_n154# VSUBS 0.05fF
C40 a_n63_n154# VSUBS 0.05fF
C41 a_n159_n154# VSUBS 0.05fF
C42 a_n255_n154# VSUBS 0.05fF
C43 w_n455_n344# VSUBS 2.96fF
.ends

.subckt inverter_cp_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_AZESM8_0 in vss in in vss out out in vss in out in vss out
+ sky130_fd_pr__nfet_01v8_AZESM8
Xsky130_fd_pr__pfet_01v8_XJXT7S_0 vss vdd in in vdd in out out in in out vdd out vdd
+ in sky130_fd_pr__pfet_01v8_XJXT7S
C0 vdd out 0.29fF
C1 out in 0.85fF
C2 vdd in 0.04fF
C3 vdd vss 5.90fF
C4 out vss 1.30fF
C5 in vss 1.82fF
.ends

.subckt pfd_cp_interface vss inverter_cp_x1_2/in vdd inverter_cp_x1_0/out Down QA
+ QB nDown Up nUp
Xinverter_cp_x2_0 nDown Down vss vdd inverter_cp_x2
Xinverter_cp_x2_1 Up nUp vss vdd inverter_cp_x2
Xtrans_gate_0 nDown vss inverter_cp_x1_0/out vdd trans_gate
Xinverter_cp_x1_0 inverter_cp_x1_0/out QB vss vdd inverter_cp_x1
Xinverter_cp_x1_2 Up inverter_cp_x1_2/in vss vdd inverter_cp_x1
Xinverter_cp_x1_1 inverter_cp_x1_2/in QA vss vdd inverter_cp_x1
C0 vdd QB 0.02fF
C1 vdd QA 0.02fF
C2 Up inverter_cp_x1_2/in 0.12fF
C3 Up nUp 0.20fF
C4 vdd Up 0.60fF
C5 Down vdd 0.09fF
C6 Down nDown 0.23fF
C7 Down inverter_cp_x1_0/out 0.12fF
C8 vdd inverter_cp_x1_2/in 0.42fF
C9 vdd nUp 0.14fF
C10 vdd nDown 0.80fF
C11 vdd inverter_cp_x1_0/out 0.25fF
C12 inverter_cp_x1_0/out nDown 0.11fF
C13 inverter_cp_x1_2/in vss 2.01fF
C14 QA vss 1.09fF
C15 inverter_cp_x1_0/out vss 2.00fF
C16 QB vss 1.09fF
C17 vdd vss 28.96fF
C18 nUp vss 1.32fF
C19 Up vss 2.53fF
C20 Down vss 1.26fF
C21 nDown vss 2.98fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4F35BC VSUBS a_n129_n90# w_n359_n309# a_n63_n116#
+ a_n159_n207# a_63_n90# a_n33_n90# a_n221_n90# a_159_n90#
X0 a_159_n90# a_n63_n116# a_63_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n129_n90# a_n159_n207# a_n221_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X2 a_63_n90# a_n159_n207# a_n33_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3 a_n33_n90# a_n63_n116# a_n129_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_n129_n90# w_n359_n309# 0.06fF
C1 a_n129_n90# a_159_n90# 0.06fF
C2 w_n359_n309# a_159_n90# 0.09fF
C3 a_63_n90# a_n129_n90# 0.09fF
C4 a_63_n90# w_n359_n309# 0.06fF
C5 a_63_n90# a_159_n90# 0.26fF
C6 a_n33_n90# a_n221_n90# 0.09fF
C7 a_n129_n90# a_n33_n90# 0.26fF
C8 a_n33_n90# w_n359_n309# 0.05fF
C9 a_n33_n90# a_159_n90# 0.09fF
C10 a_n159_n207# a_n63_n116# 0.12fF
C11 a_n129_n90# a_n221_n90# 0.26fF
C12 a_63_n90# a_n33_n90# 0.26fF
C13 a_n221_n90# w_n359_n309# 0.09fF
C14 a_n221_n90# a_159_n90# 0.04fF
C15 a_63_n90# a_n221_n90# 0.06fF
C16 a_159_n90# VSUBS 0.03fF
C17 a_63_n90# VSUBS 0.03fF
C18 a_n33_n90# VSUBS 0.03fF
C19 a_n129_n90# VSUBS 0.03fF
C20 a_n221_n90# VSUBS 0.03fF
C21 a_n159_n207# VSUBS 0.30fF
C22 a_n63_n116# VSUBS 0.37fF
C23 w_n359_n309# VSUBS 2.23fF
.ends

.subckt sky130_fd_pr__nfet_01v8_C3YG4M a_n33_n45# a_33_n71# a_n129_71# w_n263_n255#
+ a_n125_n45# a_63_n45#
X0 a_63_n45# a_33_n71# a_n33_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n129_71# a_n125_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_n33_n45# a_63_n45# 0.13fF
C1 a_n33_n45# a_n125_n45# 0.13fF
C2 a_n125_n45# a_63_n45# 0.05fF
C3 a_n129_71# a_33_n71# 0.04fF
C4 a_63_n45# w_n263_n255# 0.04fF
C5 a_n33_n45# w_n263_n255# 0.04fF
C6 a_n125_n45# w_n263_n255# 0.04fF
C7 a_33_n71# w_n263_n255# 0.11fF
C8 a_n129_71# w_n263_n255# 0.14fF
.ends

.subckt nor_pfd vdd sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss A B
Xsky130_fd_pr__pfet_01v8_4F35BC_0 vss sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vdd B A sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out vdd vdd sky130_fd_pr__pfet_01v8_4F35BC
Xsky130_fd_pr__nfet_01v8_C3YG4M_0 out B A vss vss vss sky130_fd_pr__nfet_01v8_C3YG4M
C0 out A 0.06fF
C1 B A 0.24fF
C2 vdd sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.02fF
C3 out sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.08fF
C4 vdd A 0.09fF
C5 vdd sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.02fF
C6 B out 0.40fF
C7 vdd out 0.11fF
C8 sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C9 out vss 0.45fF
C10 sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C11 A vss 0.83fF
C12 B vss 1.09fF
C13 vdd vss 3.79fF
.ends

.subckt dff_pfd vdd vss nor_pfd_2/A Q CLK nor_pfd_3/A Reset nor_pfd_2/B
Xnor_pfd_0 vdd nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_2/A nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss CLK Q nor_pfd
Xnor_pfd_1 vdd nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# Q nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss nor_pfd_2/A nor_pfd_3/A nor_pfd
Xnor_pfd_2 vdd nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_3/A nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss nor_pfd_2/A nor_pfd_2/B nor_pfd
Xnor_pfd_3 vdd nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_2/B nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss nor_pfd_3/A Reset nor_pfd
C0 Q vdd 0.08fF
C1 nor_pfd_3/A nor_pfd_2/B 0.58fF
C2 nor_pfd_2/A nor_pfd_2/B 0.05fF
C3 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vdd 0.06fF
C4 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vdd 0.06fF
C5 vdd nor_pfd_2/B 0.02fF
C6 Q Reset 0.14fF
C7 Q nor_pfd_2/B 2.22fF
C8 nor_pfd_3/A nor_pfd_2/A 0.38fF
C9 Reset nor_pfd_2/B 0.43fF
C10 Q CLK 0.04fF
C11 vdd nor_pfd_3/A 0.09fF
C12 vdd nor_pfd_2/A -0.01fF
C13 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vdd 0.06fF
C14 Q nor_pfd_3/A 0.98fF
C15 vdd nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.06fF
C16 Q nor_pfd_2/A 1.38fF
C17 vdd nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.06fF
C18 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vdd 0.06fF
C19 nor_pfd_3/A Reset 0.12fF
C20 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C21 nor_pfd_2/B vss 1.42fF
C22 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C23 nor_pfd_3/A vss 3.16fF
C24 Reset vss 1.48fF
C25 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C26 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C27 nor_pfd_2/A vss 2.56fF
C28 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C29 Q vss 2.77fF
C30 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C31 vdd vss 16.42fF
C32 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C33 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C34 CLK vss 0.95fF
.ends

.subckt sky130_fd_pr__nfet_01v8_ZCYAJJ w_n359_n255# a_n33_n45# a_n159_n173# a_n221_n45#
+ a_159_n45# a_n63_n71# a_n129_n45# a_63_n45#
X0 a_63_n45# a_n159_n173# a_n33_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n63_n71# a_n129_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X2 a_159_n45# a_n63_n71# a_63_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X3 a_n129_n45# a_n159_n173# a_n221_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_n221_n45# a_63_n45# 0.03fF
C1 a_n33_n45# a_63_n45# 0.13fF
C2 a_63_n45# a_159_n45# 0.13fF
C3 a_n33_n45# a_n221_n45# 0.05fF
C4 a_n129_n45# a_63_n45# 0.05fF
C5 a_n221_n45# a_159_n45# 0.02fF
C6 a_n129_n45# a_n221_n45# 0.13fF
C7 a_n159_n173# a_n63_n71# 0.10fF
C8 a_n33_n45# a_159_n45# 0.05fF
C9 a_n129_n45# a_n33_n45# 0.13fF
C10 a_n129_n45# a_159_n45# 0.03fF
C11 a_159_n45# w_n359_n255# 0.04fF
C12 a_63_n45# w_n359_n255# 0.05fF
C13 a_n33_n45# w_n359_n255# 0.05fF
C14 a_n129_n45# w_n359_n255# 0.05fF
C15 a_n221_n45# w_n359_n255# 0.08fF
C16 a_n159_n173# w_n359_n255# 0.31fF
C17 a_n63_n71# w_n359_n255# 0.31fF
.ends

.subckt sky130_fd_pr__pfet_01v8_7T83YG VSUBS a_n125_n90# a_63_n90# a_33_n187# a_n99_n187#
+ a_n33_n90# w_n263_n309#
X0 a_63_n90# a_33_n187# a_n33_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n33_n90# a_n99_n187# a_n125_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_n125_n90# a_63_n90# 0.09fF
C1 a_63_n90# a_n33_n90# 0.26fF
C2 a_n125_n90# a_n33_n90# 0.26fF
C3 a_n99_n187# a_33_n187# 0.04fF
C4 a_63_n90# VSUBS 0.03fF
C5 a_n33_n90# VSUBS 0.03fF
C6 a_n125_n90# VSUBS 0.03fF
C7 a_33_n187# VSUBS 0.12fF
C8 a_n99_n187# VSUBS 0.12fF
C9 w_n263_n309# VSUBS 1.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_ZXAV3F a_n73_n45# a_n33_67# a_15_n45# w_n211_n255#
X0 a_15_n45# a_n33_67# a_n73_n45# w_n211_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_n73_n45# a_15_n45# 0.16fF
C1 a_15_n45# w_n211_n255# 0.08fF
C2 a_n73_n45# w_n211_n255# 0.06fF
C3 a_n33_67# w_n211_n255# 0.10fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4F7GBC VSUBS a_n51_n187# a_n73_n90# a_15_n90# w_n211_n309#
X0 a_15_n90# a_n51_n187# a_n73_n90# w_n211_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_n73_n90# w_n211_n309# 0.04fF
C1 a_15_n90# w_n211_n309# 0.09fF
C2 a_15_n90# a_n73_n90# 0.31fF
C3 a_15_n90# VSUBS 0.03fF
C4 a_n73_n90# VSUBS 0.03fF
C5 a_n51_n187# VSUBS 0.12fF
C6 w_n211_n309# VSUBS 1.24fF
.ends

.subckt and_pfd a_656_410# vss out vdd A B
Xsky130_fd_pr__nfet_01v8_ZCYAJJ_0 vss a_656_410# A vss vss B sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45#
+ sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# sky130_fd_pr__nfet_01v8_ZCYAJJ
Xsky130_fd_pr__pfet_01v8_7T83YG_0 vss vdd vdd B A a_656_410# vdd sky130_fd_pr__pfet_01v8_7T83YG
Xsky130_fd_pr__nfet_01v8_ZXAV3F_0 vss a_656_410# out vss sky130_fd_pr__nfet_01v8_ZXAV3F
Xsky130_fd_pr__pfet_01v8_4F7GBC_0 vss a_656_410# vdd out vdd sky130_fd_pr__pfet_01v8_4F7GBC
C0 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# out 0.03fF
C1 A vdd 0.05fF
C2 a_656_410# B 0.30fF
C3 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# a_656_410# 0.07fF
C4 a_656_410# out 0.20fF
C5 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# B 0.02fF
C6 out vdd 0.10fF
C7 A B 0.33fF
C8 a_656_410# vdd 0.20fF
C9 A a_656_410# 0.04fF
C10 vdd vss 4.85fF
C11 out vss 0.47fF
C12 a_656_410# vss 1.00fF
C13 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.13fF
C14 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.10fF
C15 A vss 0.85fF
C16 B vss 0.95fF
.ends

.subckt PFD vss vdd Reset Down Up A B
Xdff_pfd_0 vdd vss dff_pfd_0/nor_pfd_2/A Up A dff_pfd_0/nor_pfd_3/A Reset dff_pfd_0/nor_pfd_2/B
+ dff_pfd
Xdff_pfd_1 vdd vss dff_pfd_1/nor_pfd_2/A Down B dff_pfd_1/nor_pfd_3/A Reset dff_pfd_1/nor_pfd_2/B
+ dff_pfd
Xand_pfd_0 and_pfd_0/a_656_410# vss Reset vdd Up Down and_pfd
C0 vdd dff_pfd_1/nor_pfd_3/A 0.08fF
C1 vdd Down 0.08fF
C2 Down Up 0.06fF
C3 vdd dff_pfd_1/nor_pfd_2/B 0.04fF
C4 vdd dff_pfd_0/nor_pfd_3/A 0.08fF
C5 vdd dff_pfd_0/nor_pfd_2/B 0.11fF
C6 vdd Reset 0.02fF
C7 vdd dff_pfd_0/nor_pfd_2/A 0.13fF
C8 vdd Up 1.62fF
C9 vdd dff_pfd_1/nor_pfd_2/A 0.13fF
C10 and_pfd_0/a_656_410# vss 0.99fF
C11 and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C12 and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.05fF
C13 dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C14 dff_pfd_1/nor_pfd_2/B vss 1.51fF
C15 dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C16 dff_pfd_1/nor_pfd_3/A vss 3.14fF
C17 dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C18 dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C19 dff_pfd_1/nor_pfd_2/A vss 2.56fF
C20 dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C21 Down vss 3.74fF
C22 dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C23 vdd vss 44.73fF
C24 dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C25 dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C26 B vss 1.07fF
C27 dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C28 dff_pfd_0/nor_pfd_2/B vss 1.40fF
C29 dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C30 dff_pfd_0/nor_pfd_3/A vss 3.14fF
C31 Reset vss 3.85fF
C32 dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C33 dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C34 dff_pfd_0/nor_pfd_2/A vss 2.56fF
C35 dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C36 Up vss 3.18fF
C37 dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C38 dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C39 dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C40 A vss 1.07fF
.ends

.subckt top_pll_v3 clk_d vdd s_0 charge_pump_0/w_2544_775# out_by_2 s_0_n in_ref ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd
+ buffer_salida_0/a_3996_n100# vss vco_vctrl s_1 ring_osc_0/csvco_branch_2/vbp lf_vc
+ vco_D0 lf_D0 buffer_salida_0/a_678_n100# ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd
+ loop_filter_v2_0/cap3_loop_filter_0/in charge_pump_0/w_1008_774# iref_cp ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd
+ Down out_to_div clk_1 out_div nDown s_1_n out_to_pad MC Up clk_0 freq_div_0/prescaler_23_0/nCLK_23
+ biasp nUp n_clk_0
Xcharge_pump_0 vss pswitch nswitch vco_vctrl vdd biasp nUp Down charge_pump_0/w_2544_775#
+ iref_cp nDown Up charge_pump_0/w_1008_774# vss charge_pump
Xdiv_by_2_0 vss vdd n_out_div_2 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in out_by_2
+ n_out_by_2 out_buffer_div_2 out_to_div out_div_2 n_out_buffer_div_2 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_2
Xloop_filter_v2_0 lf_vc lf_D0 vco_vctrl vss loop_filter_v2_0/cap3_loop_filter_0/in
+ loop_filter_v2
Xbuffer_salida_0 buffer_salida_0/a_678_n100# buffer_salida_0/a_3996_n100# out_to_pad
+ vdd out_to_buffer vss buffer_salida
Xfreq_div_0 clk_0 vss out_by_2 n_clk_0 vdd freq_div_0/prescaler_23_0/Q2 s_0 s_1_n
+ s_1 freq_div_0/prescaler_23_0/nCLK_23 MC clk_d freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280#
+ s_0_n clk_pre freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/D
+ freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/nD clk_1 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280#
+ clk_out_mux21 n_clk_1 out_div freq_div_0/div_by_5_0/Q1 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D
+ freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD
+ clk_2_f n_out_by_2 clk_5 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/nD freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D
+ freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/D freq_div
Xring_osc_0 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vco_vctrl vss ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd
+ ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vdd ring_osc_0/csvco_branch_2/vbp
+ ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vco_D0 ring_osc_0/csvco_branch_2/cap_vco_0/t
+ vco_out ring_osc
Xring_osc_buffer_0 vss vco_out vdd out_first_buffer out_to_div out_to_buffer ring_osc_buffer
Xpfd_cp_interface_0 vss pfd_cp_interface_0/inverter_cp_x1_2/in vdd pfd_cp_interface_0/inverter_cp_x1_0/out
+ Down QA QB nDown Up nUp pfd_cp_interface
XPFD_0 vss vdd pfd_reset QB QA in_ref out_div PFD
C0 pswitch nDown 0.53fF
C1 nDown nUp -0.09fF
C2 vco_vctrl freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/D 0.53fF
C3 vco_vctrl freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/nD 1.23fF
C4 charge_pump_0/w_2544_775# nDown 0.05fF
C5 s_1_n out_div 0.10fF
C6 vco_vctrl freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D 0.65fF
C7 vdd QA -0.04fF
C8 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vco_vctrl 0.82fF
C9 pswitch Up 1.98fF
C10 Up nUp 2.72fF
C11 vco_vctrl freq_div_0/prescaler_23_0/nCLK_23 0.06fF
C12 vdd clk_0 0.13fF
C13 vdd ring_osc_0/csvco_branch_2/vbp 0.03fF
C14 vdd nDown 0.22fF
C15 s_0_n n_out_by_2 0.14fF
C16 vco_vctrl n_clk_1 0.23fF
C17 clk_d out_div 0.64fF
C18 s_0 out_to_div 0.94fF
C19 pswitch nUp 0.93fF
C20 vco_D0 vdd 0.03fF
C21 clk_1 n_out_by_2 -0.10fF
C22 nswitch nDown 0.76fF
C23 lf_vc MC 0.20fF
C24 vco_vctrl clk_0 -0.26fF
C25 vco_vctrl ring_osc_0/csvco_branch_2/vbp 0.26fF
C26 vdd Up 0.28fF
C27 out_div s_1 0.37fF
C28 vco_vctrl ring_osc_0/csvco_branch_0/inverter_csvco_0/vss 0.04fF
C29 s_0 n_out_by_2 0.14fF
C30 out_to_div out_to_buffer 0.13fF
C31 iref_cp Down 0.09fF
C32 biasp Down 1.24fF
C33 nDown Down 2.55fF
C34 vdd nUp 0.05fF
C35 vdd ring_osc_0/csvco_branch_2/cap_vco_0/t 0.02fF
C36 ring_osc_0/csvco_branch_2/cap_vco_0/t out_first_buffer 0.03fF
C37 vco_vctrl MC 0.33fF
C38 vco_vctrl freq_div_0/div_by_5_0/Q1 0.10fF
C39 vco_vctrl freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/D 0.09fF
C40 buffer_salida_0/a_678_n100# vdd 0.24fF
C41 vco_vctrl freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD -0.42fF
C42 charge_pump_0/w_2544_775# Down -0.23fF
C43 vco_vctrl s_0_n 0.34fF
C44 vco_vctrl vdd 0.82fF
C45 vco_vctrl clk_1 -0.04fF
C46 biasp nDown 0.26fF
C47 vdd pfd_cp_interface_0/inverter_cp_x1_2/in 0.01fF
C48 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D vco_vctrl -0.42fF
C49 buffer_salida_0/a_678_n100# out_to_buffer 0.21fF
C50 vdd out_to_buffer 0.07fF
C51 vco_vctrl s_0 0.45fF
C52 nswitch Down 0.54fF
C53 biasp Up 0.26fF
C54 vco_vctrl freq_div_0/prescaler_23_0/Q2 0.06fF
C55 vco_vctrl freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD 0.15fF
C56 vco_vctrl freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# 0.34fF
C57 vco_vctrl freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/nD 0.09fF
C58 out_by_2 n_out_by_2 0.27fF
C59 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# vco_vctrl 0.17fF
C60 biasp nUp -0.16fF
C61 PFD_0/and_pfd_0/a_656_410# vss 0.96fF
C62 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C63 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.07fF
C64 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C65 PFD_0/dff_pfd_1/nor_pfd_2/B vss 1.40fF
C66 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C67 PFD_0/dff_pfd_1/nor_pfd_3/A vss 3.14fF
C68 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C69 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C70 PFD_0/dff_pfd_1/nor_pfd_2/A vss 2.55fF
C71 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C72 QB vss 3.15fF
C73 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C74 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C75 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C76 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C77 PFD_0/dff_pfd_0/nor_pfd_2/B vss 1.40fF
C78 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C79 PFD_0/dff_pfd_0/nor_pfd_3/A vss 3.14fF
C80 pfd_reset vss 1.87fF
C81 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C82 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C83 PFD_0/dff_pfd_0/nor_pfd_2/A vss 2.55fF
C84 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C85 QA vss 3.49fF
C86 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C87 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C88 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C89 in_ref vss 0.84fF
C90 pfd_cp_interface_0/inverter_cp_x1_2/in vss 1.85fF
C91 pfd_cp_interface_0/inverter_cp_x1_0/out vss 1.87fF
C92 nUp vss 0.12fF
C93 Up vss -4.26fF
C94 Down vss 1.89fF
C95 nDown vss 2.80fF
C96 out_first_buffer vss 2.15fF
C97 out_to_buffer vss 1.92fF
C98 out_to_div vss 8.72fF
C99 ring_osc_0/csvco_branch_2/in vss 1.60fF
C100 ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C101 ring_osc_0/csvco_branch_1/cap_vco_0/t vss 7.10fF
C102 ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vss 0.52fF
C103 ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C104 ring_osc_0/csvco_branch_2/cap_vco_0/t vss 7.10fF
C105 ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vss 0.52fF
C106 ring_osc_0/csvco_branch_1/in vss 1.58fF
C107 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C108 vco_out vss 1.65fF
C109 vco_D0 vss -4.72fF
C110 ring_osc_0/csvco_branch_0/cap_vco_0/t vss 7.10fF
C111 ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vss 0.52fF
C112 ring_osc_0/csvco_branch_2/vbp vss 0.38fF
C113 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_1/a_63_368# vss 0.37fF
C114 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C115 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_0/X vss 0.49fF
C116 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C117 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C118 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C119 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C120 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C121 freq_div_0/prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C122 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C123 freq_div_0/prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C124 freq_div_0/prescaler_23_0/DFlipFlop_1/D vss 1.90fF
C125 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C126 freq_div_0/prescaler_23_0/Q2_d vss -0.69fF
C127 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C128 freq_div_0/prescaler_23_0/DFlipFlop_2/nQ vss 0.48fF
C129 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C130 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C131 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C132 freq_div_0/prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C133 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C134 freq_div_0/prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C135 freq_div_0/prescaler_23_0/Q2 vss 0.55fF
C136 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C137 freq_div_0/prescaler_23_0/Q1 vss 0.07fF
C138 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C139 n_clk_0 vss -7.01fF
C140 freq_div_0/prescaler_23_0/DFlipFlop_0/nQ vss 0.48fF
C141 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C142 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C143 clk_0 vss -0.37fF
C144 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C145 freq_div_0/prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C146 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C147 freq_div_0/prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C148 freq_div_0/prescaler_23_0/nCLK_23 vss -1.02fF
C149 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C150 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_1/X vss -1.01fF
C151 MC vss -1.42fF
C152 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_304_74# vss 0.36fF
C153 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_27_112# vss 0.65fF
C154 n_out_by_2 vss 4.87fF
C155 s_0_n vss -4.09fF
C156 out_by_2 vss 4.52fF
C157 s_0 vss 5.50fF
C158 freq_div_0/div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C159 freq_div_0/div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.38fF
C160 freq_div_0/div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C161 freq_div_0/div_by_5_0/Q1_shift vss -0.36fF
C162 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.57fF
C163 freq_div_0/div_by_5_0/DFlipFlop_3/nQ vss 0.48fF
C164 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_1/D vss -1.73fF
C165 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C166 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C167 freq_div_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C168 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_0/D vss 0.96fF
C169 freq_div_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C170 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C171 freq_div_0/div_by_5_0/Q1 vss 4.35fF
C172 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C173 freq_div_0/div_by_5_0/DFlipFlop_2/nQ vss 0.48fF
C174 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C175 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C176 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C177 freq_div_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C178 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C179 freq_div_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C180 freq_div_0/div_by_5_0/DFlipFlop_2/D vss 3.13fF
C181 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C182 freq_div_0/div_by_5_0/Q0 vss 0.29fF
C183 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C184 freq_div_0/div_by_5_0/nQ0 vss 0.99fF
C185 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C186 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C187 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C188 freq_div_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C189 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C190 freq_div_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C191 freq_div_0/div_by_5_0/DFlipFlop_1/D vss 3.64fF
C192 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C193 freq_div_0/div_by_5_0/DFlipFlop_0/Q vss -0.94fF
C194 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C195 n_clk_1 vss -0.56fF
C196 freq_div_0/div_by_5_0/nQ2 vss 1.38fF
C197 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C198 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C199 clk_1 vss -2.21fF
C200 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C201 freq_div_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C202 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C203 freq_div_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C204 freq_div_0/div_by_5_0/DFlipFlop_0/D vss 3.96fF
C205 vdd vss 587.93fF
C206 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C207 freq_div_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C208 freq_div_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.40fF
C209 s_1_n vss -2.04fF
C210 out_div vss 3.70fF
C211 clk_d vss 1.27fF
C212 s_1 vss 1.72fF
C213 freq_div_0/inverter_min_x4_0/in vss 2.71fF
C214 clk_5 vss -0.22fF
C215 clk_out_mux21 vss 3.89fF
C216 clk_pre vss 1.69fF
C217 freq_div_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C218 freq_div_0/div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C219 freq_div_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C220 freq_div_0/div_by_2_0/DFlipFlop_0/nCLK vss 1.03fF
C221 clk_2_f vss 3.30fF
C222 freq_div_0/div_by_2_0/o1 vss 2.08fF
C223 freq_div_0/div_by_2_0/nCLK_2 vss 1.04fF
C224 freq_div_0/div_by_2_0/o2 vss 2.08fF
C225 freq_div_0/div_by_2_0/out_div vss -0.82fF
C226 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C227 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C228 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C229 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C230 freq_div_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C231 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C232 freq_div_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C233 freq_div_0/div_by_2_0/nout_div vss 2.62fF
C234 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C235 out_to_pad vss 7.15fF
C236 buffer_salida_0/a_3996_n100# vss 48.29fF
C237 buffer_salida_0/a_678_n100# vss 13.38fF
C238 lf_vc vss -60.88fF
C239 loop_filter_v2_0/res_loop_filter_2/out vss 7.90fF
C240 lf_D0 vss 0.01fF
C241 loop_filter_v2_0/cap3_loop_filter_0/in vss -12.03fF
C242 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C243 div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C244 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C245 div_by_2_0/DFlipFlop_0/nCLK vss 1.03fF
C246 out_buffer_div_2 vss 1.57fF
C247 n_out_buffer_div_2 vss 1.57fF
C248 out_div_2 vss -0.70fF
C249 div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C250 div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C251 div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C252 div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C253 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C254 div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C255 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C256 n_out_div_2 vss 2.11fF
C257 div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C258 nswitch vss 4.61fF
C259 biasp vss 5.46fF
C260 iref_cp vss 2.44fF
C261 vco_vctrl vss -30.24fF
C262 pswitch vss 2.72fF
.ends

.subckt loop_filter vc_pex in vss
Xcap1_loop_filter_0 vss vc_pex vss cap1_loop_filter
Xcap2_loop_filter_0 vss in vss cap2_loop_filter
Xres_loop_filter_0 vss res_loop_filter_2/out in res_loop_filter
Xres_loop_filter_1 vss res_loop_filter_2/out vc_pex res_loop_filter
Xres_loop_filter_2 vss res_loop_filter_2/out vc_pex res_loop_filter
C0 in vc_pex 0.18fF
C1 vc_pex vss -38.13fF
C2 res_loop_filter_2/out vss 8.49fF
C3 in vss -18.79fF
.ends

.subckt top_pll_v1 vco_vctrl ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vdd charge_pump_0/w_2544_775#
+ pswitch biasp ring_osc_0/csvco_branch_2/vbp in_ref Down w_13905_n238# vss vco_D0
+ QA ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd iref_cp out_to_div nDown out_to_pad
+ ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd Up nUp
Xloop_filter_0 lf_vc vco_vctrl vss loop_filter
Xcharge_pump_0 vss pswitch nswitch vco_vctrl vdd biasp nUp Down charge_pump_0/w_2544_775#
+ iref_cp nDown Up charge_pump_0/w_1008_774# charge_pump_0/w_6648_570# charge_pump
Xdiv_by_2_0 vss vdd n_out_div_2 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in out_by_2
+ n_out_by_2 out_buffer_div_2 out_to_div out_div_2 n_out_buffer_div_2 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_2
Xbuffer_salida_0 buffer_salida_0/a_678_n100# buffer_salida_0/a_3996_n100# out_to_pad
+ vdd out_to_buffer vss buffer_salida
Xring_osc_0 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vco_vctrl vss ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd
+ ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vdd ring_osc_0/csvco_branch_2/vbp
+ ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vco_D0 ring_osc_0/csvco_branch_2/cap_vco_0/t
+ vco_out ring_osc
Xring_osc_buffer_0 vss vco_out vdd out_first_buffer out_to_div out_to_buffer ring_osc_buffer
Xdiv_by_5_0 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in n_out_by_2
+ div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/DFlipFlop_0/latch_diff_1/nD
+ vss vdd div_by_5_0/DFlipFlop_2/latch_diff_0/nD div_5_Q0 div_5_Q1 out_by_2 div_by_5_0/DFlipFlop_0/Q
+ div_by_5_0/DFlipFlop_2/latch_diff_1/D div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# div_5_nQ0 div_by_5_0/DFlipFlop_3/latch_diff_0/D
+ div_by_5_0/DFlipFlop_3/latch_diff_1/nD div_by_5_0/DFlipFlop_1/latch_diff_1/nD div_by_5_0/DFlipFlop_1/latch_diff_0/nD
+ div_by_5_0/DFlipFlop_1/latch_diff_0/D div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280#
+ out_div_by_5 div_5_Q1_shift div_5_nQ2 div_by_5_0/DFlipFlop_2/D div_by_5_0/DFlipFlop_2/latch_diff_1/nD
+ div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out div_by_5_0/DFlipFlop_1/latch_diff_1/D
+ div_by_5_0/DFlipFlop_1/D div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ div_by_5_0/DFlipFlop_0/latch_diff_0/nD div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368#
+ div_by_5_0/DFlipFlop_0/D div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_0/latch_diff_1/D div_by_5_0/DFlipFlop_2/nQ div_by_5_0/DFlipFlop_3/latch_diff_0/nD
+ div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out div_by_5_0/DFlipFlop_2/latch_diff_0/D
+ div_by_5_0/DFlipFlop_0/latch_diff_0/D div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ div_by_5_0/DFlipFlop_3/latch_diff_1/D div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368#
+ div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136#
+ div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_152_368# div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# div_by_5_0/DFlipFlop_3/nQ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136#
+ div_by_5
Xpfd_cp_interface_0 vss pfd_cp_interface_0/inverter_cp_x1_2/in vdd pfd_cp_interface_0/inverter_cp_x1_0/out
+ Down QA QB nDown Up nUp pfd_cp_interface
XPFD_0 vss vdd pfd_reset QB QA in_ref out_div_by_5 PFD
C0 div_5_nQ2 n_out_by_2 0.10fF
C1 vdd pfd_cp_interface_0/inverter_cp_x1_2/in 0.01fF
C2 div_5_nQ2 out_by_2 0.16fF
C3 lf_vc vdd 0.02fF
C4 div_by_5_0/DFlipFlop_0/latch_diff_0/D n_out_by_2 0.24fF
C5 nDown biasp 0.26fF
C6 out_by_2 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.28fF
C7 vdd out_to_buffer 0.07fF
C8 vdd nUp 0.05fF
C9 n_out_by_2 div_by_5_0/DFlipFlop_0/Q -0.23fF
C10 Down iref_cp 0.09fF
C11 n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/D 0.17fF
C12 out_by_2 div_by_5_0/DFlipFlop_0/Q 0.09fF
C13 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in out_to_div -0.16fF
C14 out_to_div vdd 0.21fF
C15 biasp Down 1.24fF
C16 n_out_by_2 div_by_5_0/DFlipFlop_1/D 0.22fF
C17 out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/D 0.33fF
C18 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in n_out_by_2 -0.51fF
C19 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# 0.02fF
C20 nDown Down 2.55fF
C21 out_by_2 div_by_5_0/DFlipFlop_1/D 0.38fF
C22 out_by_2 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# 0.10fF
C23 div_by_5_0/DFlipFlop_3/latch_diff_1/nD n_out_by_2 0.10fF
C24 buffer_salida_0/a_678_n100# vdd 0.24fF
C25 out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/nD 0.23fF
C26 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392# n_out_by_2 0.01fF
C27 n_out_by_2 div_5_Q0 -0.12fF
C28 vdd Up 0.28fF
C29 out_div_by_5 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# 0.18fF
C30 n_out_by_2 div_5_Q1 1.04fF
C31 pswitch nUp 0.85fF
C32 out_by_2 div_5_Q0 0.09fF
C33 out_by_2 div_5_Q1 0.42fF
C34 out_div_by_5 div_5_Q1_shift 0.05fF
C35 out_to_div out_to_buffer 0.13fF
C36 n_out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_0/nD 0.11fF
C37 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# vco_vctrl -0.11fF
C38 n_out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_0/D 0.12fF
C39 n_out_by_2 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.27fF
C40 buffer_salida_0/a_678_n100# out_to_buffer 0.22fF
C41 n_out_by_2 div_by_5_0/DFlipFlop_0/D -1.48fF
C42 n_out_by_2 div_by_5_0/DFlipFlop_2/nQ 0.10fF
C43 n_out_by_2 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out -0.11fF
C44 vdd iref_cp 0.15fF
C45 out_by_2 div_by_5_0/DFlipFlop_0/D 0.35fF
C46 div_5_Q0 vco_vctrl 0.48fF
C47 n_out_by_2 div_by_5_0/DFlipFlop_2/D 0.19fF
C48 pswitch Up 1.98fF
C49 out_by_2 div_by_5_0/DFlipFlop_2/nQ 0.23fF
C50 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# 0.12fF
C51 ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vco_vctrl 0.04fF
C52 n_out_by_2 vco_vctrl 0.52fF
C53 vco_vctrl div_5_Q1 0.14fF
C54 Up nUp 2.72fF
C55 out_by_2 div_by_5_0/DFlipFlop_2/D 0.22fF
C56 n_out_by_2 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in -0.20fF
C57 nDown vdd 0.22fF
C58 out_by_2 vco_vctrl 0.53fF
C59 div_5_nQ0 n_out_by_2 0.10fF
C60 vco_D0 vdd 0.03fF
C61 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136# out_by_2 -0.02fF
C62 div_5_nQ0 out_by_2 0.32fF
C63 out_by_2 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out -0.04fF
C64 n_out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/nD 0.24fF
C65 n_out_by_2 vdd 1.03fF
C66 out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/nD 0.09fF
C67 n_out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/D 0.24fF
C68 out_by_2 vdd 0.97fF
C69 vco_vctrl div_by_5_0/DFlipFlop_0/D -0.45fF
C70 nDown nswitch 0.76fF
C71 out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_0/nD 0.17fF
C72 out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/D 0.09fF
C73 vdd ring_osc_0/csvco_branch_2/cap_vco_0/t 0.02fF
C74 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vco_vctrl -0.36fF
C75 vco_vctrl ring_osc_0/csvco_branch_2/vbp 0.26fF
C76 out_div_by_5 div_5_Q1 0.01fF
C77 out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_0/nD 0.10fF
C78 biasp nUp -0.17fF
C79 nDown pswitch 0.53fF
C80 n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.33fF
C81 out_first_buffer ring_osc_0/csvco_branch_2/cap_vco_0/t 0.03fF
C82 Down nswitch 0.54fF
C83 nDown nUp -0.09fF
C84 out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.17fF
C85 n_out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_1/nD 0.24fF
C86 out_by_2 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out 0.09fF
C87 vdd div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out 0.04fF
C88 out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_1/nD 0.09fF
C89 vdd div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# 0.03fF
C90 vdd ring_osc_0/csvco_branch_2/vbp 0.03fF
C91 vdd vco_vctrl -1.02fF
C92 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# 0.03fF
C93 biasp Up 0.26fF
C94 n_out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_0/D 0.12fF
C95 n_out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_1/D 0.10fF
C96 vco_vctrl nswitch -0.06fF
C97 out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_1/D 0.23fF
C98 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# -0.05fF
C99 n_out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/D 0.10fF
C100 out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_0/nD 0.10fF
C101 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out out_to_div -0.12fF
C102 out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/D 0.23fF
C103 out_div_by_5 vdd 0.28fF
C104 nUp vco_vctrl 0.02fF
C105 QA vdd -0.04fF
C106 div_by_5_0/DFlipFlop_3/latch_diff_0/D out_by_2 0.11fF
C107 out_by_2 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in -0.22fF
C108 PFD_0/and_pfd_0/a_656_410# vss 0.96fF
C109 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C110 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.07fF
C111 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C112 PFD_0/dff_pfd_1/nor_pfd_2/B vss 1.40fF
C113 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C114 PFD_0/dff_pfd_1/nor_pfd_3/A vss 3.14fF
C115 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C116 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C117 PFD_0/dff_pfd_1/nor_pfd_2/A vss 2.55fF
C118 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C119 QB vss 4.46fF
C120 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C121 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C122 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C123 out_div_by_5 vss -0.40fF
C124 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C125 PFD_0/dff_pfd_0/nor_pfd_2/B vss 1.40fF
C126 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C127 PFD_0/dff_pfd_0/nor_pfd_3/A vss 3.14fF
C128 pfd_reset vss 2.17fF
C129 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C130 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C131 PFD_0/dff_pfd_0/nor_pfd_2/A vss 2.55fF
C132 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C133 QA vss 4.31fF
C134 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C135 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C136 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C137 in_ref vss 1.19fF
C138 pfd_cp_interface_0/inverter_cp_x1_2/in vss 1.85fF
C139 pfd_cp_interface_0/inverter_cp_x1_0/out vss 1.87fF
C140 nUp vss 5.50fF
C141 Up vss 2.37fF
C142 Down vss 7.92fF
C143 nDown vss -2.20fF
C144 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C145 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.38fF
C146 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.41fF
C147 div_5_Q1_shift vss -0.14fF
C148 div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.57fF
C149 div_by_5_0/DFlipFlop_3/nQ vss 0.48fF
C150 div_by_5_0/DFlipFlop_3/latch_diff_1/D vss -1.73fF
C151 div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C152 div_by_5_0/DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C153 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C154 div_by_5_0/DFlipFlop_3/latch_diff_0/D vss 0.96fF
C155 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C156 div_by_5_0/DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C157 div_5_Q1 vss 4.28fF
C158 div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C159 div_by_5_0/DFlipFlop_2/nQ vss 0.48fF
C160 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C161 div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C162 div_by_5_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C163 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C164 div_by_5_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C165 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C166 div_by_5_0/DFlipFlop_2/D vss 3.13fF
C167 div_by_5_0/DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C168 div_5_Q0 vss 0.01fF
C169 div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C170 div_5_nQ0 vss 0.59fF
C171 div_by_5_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C172 div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C173 div_by_5_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C174 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C175 div_by_5_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C176 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C177 div_by_5_0/DFlipFlop_1/D vss 3.64fF
C178 div_by_5_0/DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C179 div_by_5_0/DFlipFlop_0/Q vss -0.94fF
C180 div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C181 n_out_by_2 vss -2.62fF
C182 div_5_nQ2 vss 1.24fF
C183 div_by_5_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C184 div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C185 out_by_2 vss -4.51fF
C186 div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C187 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C188 div_by_5_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C189 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C190 div_by_5_0/DFlipFlop_0/D vss 3.96fF
C191 vdd vss 366.82fF
C192 div_by_5_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C193 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C194 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.40fF
C195 out_first_buffer vss 2.88fF
C196 out_to_buffer vss 1.57fF
C197 out_to_div vss 4.46fF
C198 ring_osc_0/csvco_branch_2/in vss 1.60fF
C199 ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C200 ring_osc_0/csvco_branch_1/cap_vco_0/t vss 7.10fF
C201 ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vss 0.52fF
C202 ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C203 ring_osc_0/csvco_branch_2/cap_vco_0/t vss 7.10fF
C204 ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vss 0.52fF
C205 ring_osc_0/csvco_branch_1/in vss 1.58fF
C206 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C207 vco_out vss 1.01fF
C208 vco_D0 vss -4.63fF
C209 ring_osc_0/csvco_branch_0/cap_vco_0/t vss 7.10fF
C210 ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vss 0.52fF
C211 ring_osc_0/csvco_branch_2/vbp vss 0.38fF
C212 out_to_pad vss 7.50fF
C213 buffer_salida_0/a_3996_n100# vss 48.29fF
C214 buffer_salida_0/a_678_n100# vss 13.38fF
C215 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C216 div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C217 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.89fF
C218 div_by_2_0/DFlipFlop_0/nCLK vss 1.03fF
C219 out_buffer_div_2 vss 1.60fF
C220 n_out_buffer_div_2 vss 1.63fF
C221 out_div_2 vss -1.30fF
C222 div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C223 div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C224 div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C225 div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C226 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C227 div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C228 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C229 n_out_div_2 vss 1.95fF
C230 div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C231 nswitch vss 3.73fF
C232 biasp vss 5.44fF
C233 iref_cp vss 2.81fF
C234 vco_vctrl vss -19.28fF
C235 pswitch vss 3.57fF
C236 lf_vc vss -59.89fF
C237 loop_filter_0/res_loop_filter_2/out vss 7.90fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_2Y8F6P VSUBS c2_n3251_n3000# m4_n3351_n3100#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
C0 c2_n3251_n3000# m4_n3351_n3100# 72.82fF
C1 m4_n3351_n3100# VSUBS 14.58fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_8P223X VSUBS a_n2017_n1317# a_n1731_n1219# a_n1879_n1219#
+ a_n2017_n61# w_n2018_n202#
X0 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X1 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X2 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X3 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X4 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X5 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X6 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X7 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X8 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X9 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X10 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X11 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X12 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X13 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X14 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X15 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X16 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X17 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X18 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X19 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X20 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X21 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X22 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X23 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X24 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X25 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X26 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X27 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X28 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X29 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X30 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X31 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X32 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X33 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X34 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X35 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X36 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X37 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X38 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X39 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X40 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X41 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X42 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X43 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X44 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X45 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X46 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X47 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X48 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X49 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
C0 a_n2017_n61# a_n2017_n1317# 2.88fF
C1 a_n1879_n1219# w_n2018_n202# 0.25fF
C2 a_n1731_n1219# a_n1879_n1219# 19.29fF
C3 w_n2018_n202# a_n2017_n1317# 0.16fF
C4 a_n1731_n1219# a_n2017_n1317# 4.73fF
C5 a_n2017_n61# w_n2018_n202# 1.37fF
C6 a_n2017_n61# a_n1731_n1219# 5.23fF
C7 a_n1879_n1219# a_n2017_n1317# 2.66fF
C8 a_n1731_n1219# w_n2018_n202# 19.90fF
C9 a_n2017_n61# a_n1879_n1219# 0.16fF
C10 a_n1879_n1219# VSUBS 1.53fF
C11 a_n2017_n1317# VSUBS 5.03fF
C12 a_n1731_n1219# VSUBS 2.60fF
C13 a_n2017_n61# VSUBS 5.10fF
C14 w_n2018_n202# VSUBS 37.43fF
.ends

.subckt bias VSUBS vdd iref_0 iref_1 iref_2 iref_5 iref_6 iref_7 iref_8 iref_9 iref
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_5 VSUBS iref m1_20168_984# iref m1_20168_984#
+ vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_6 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_6/a_n1731_n1219#
+ iref_5 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_7 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219#
+ iref_6 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_9 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219#
+ iref_8 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_8 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219#
+ iref_7 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_10 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219#
+ iref_9 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_0 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_0/a_n1731_n1219#
+ iref_0 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_1 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219#
+ iref_1 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_2 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219#
+ iref_2 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_3 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219#
+ iref_3 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_4 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219#
+ iref_4 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
C0 m1_20168_984# sky130_fd_pr__pfet_01v8_lvt_8P223X_6/a_n1731_n1219# 0.54fF
C1 sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# iref_2 0.24fF
C2 m1_20168_984# vdd 0.25fF
C3 sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219# vdd 0.24fF
C4 sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# sky130_fd_pr__pfet_01v8_lvt_8P223X_0/a_n1731_n1219# 0.67fF
C5 sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# m1_20168_984# -0.39fF
C6 iref m1_20168_984# 0.07fF
C7 sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219# iref_6 0.24fF
C8 iref_4 iref 0.30fF
C9 sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# m1_20168_984# 0.01fF
C10 iref_4 iref_3 0.05fF
C11 iref_2 iref -0.01fF
C12 iref_9 iref_8 0.05fF
C13 iref_9 iref -0.01fF
C14 iref_2 iref_3 0.05fF
C15 sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# vdd 0.24fF
C16 iref_8 iref_7 0.05fF
C17 sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219# vdd 0.24fF
C18 iref_6 iref_7 0.05fF
C19 iref_2 iref_1 0.05fF
C20 sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219# vdd 0.24fF
C21 sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219# iref_1 0.24fF
C22 iref vdd -0.07fF
C23 iref_8 iref -0.03fF
C24 sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# iref -0.15fF
C25 iref_7 sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219# 0.24fF
C26 iref_5 sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219# 0.24fF
C27 sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# vdd 0.24fF
C28 iref_0 iref_1 0.05fF
C29 sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# iref 0.02fF
C30 iref_1 iref -0.02fF
C31 iref_5 iref_6 0.05fF
C32 iref_5 iref 0.05fF
C33 sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219# vdd 0.24fF
C34 sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219# iref_8 0.24fF
C35 sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# m1_20168_984# 0.01fF
C36 sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# iref_3 0.24fF
C37 sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219# vdd 0.24fF
C38 iref_4 VSUBS 1.17fF
C39 sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# VSUBS 2.60fF
C40 iref_3 VSUBS 0.64fF
C41 sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# VSUBS 2.60fF
C42 iref_2 VSUBS -1.26fF
C43 sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219# VSUBS 2.60fF
C44 iref_1 VSUBS -0.80fF
C45 sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# VSUBS 2.60fF
C46 iref_0 VSUBS 1.88fF
C47 iref VSUBS 32.42fF
C48 sky130_fd_pr__pfet_01v8_lvt_8P223X_0/a_n1731_n1219# VSUBS 2.60fF
C49 m1_20168_984# VSUBS 56.92fF
C50 vdd VSUBS 416.01fF
C51 iref_9 VSUBS -1.13fF
C52 sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219# VSUBS 2.60fF
C53 iref_7 VSUBS -1.38fF
C54 sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219# VSUBS 2.60fF
C55 iref_8 VSUBS -1.19fF
C56 sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219# VSUBS 2.60fF
C57 iref_6 VSUBS -1.00fF
C58 sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219# VSUBS 2.60fF
C59 iref_5 VSUBS 1.40fF
C60 sky130_fd_pr__pfet_01v8_lvt_8P223X_6/a_n1731_n1219# VSUBS 2.60fF
.ends

.subckt mimcap_decoup_1x5 VSUBS t b
Xdecap[0] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[1] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[2] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[3] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[4] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
C0 b VSUBS 68.24fF
.ends

.subckt top_pll_v2 ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd pswitch vdd charge_pump_0/w_2544_775#
+ ring_osc_0/csvco_branch_2/vbp ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd in_ref
+ vco_vctrl Down w_13905_n238# vss D0_vco iref_cp ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd
+ out_to_div DO_cap nDown biasp out_to_pad Up nUp
Xcharge_pump_0 vss pswitch nswitch vco_vctrl vdd biasp nUp Down charge_pump_0/w_2544_775#
+ iref_cp nDown Up charge_pump_0/w_1008_774# charge_pump_0/w_6648_570# charge_pump
Xdiv_by_2_0 vss vdd n_out_div_2 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in out_by_2
+ n_out_by_2 out_buffer_div_2 out_to_div out_div_2 n_out_buffer_div_2 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_2
Xloop_filter_v2_0 lf_vc DO_cap vco_vctrl vss loop_filter_v2_0/cap3_loop_filter_0/in
+ loop_filter_v2
Xbuffer_salida_0 buffer_salida_0/a_678_n100# buffer_salida_0/a_3996_n100# out_to_pad
+ vdd out_to_buffer vss buffer_salida
Xring_osc_0 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vco_vctrl vss ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd
+ ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vdd ring_osc_0/csvco_branch_2/vbp
+ ring_osc_0/csvco_branch_0/inverter_csvco_0/vss D0_vco ring_osc_0/csvco_branch_2/cap_vco_0/t
+ vco_out ring_osc
Xring_osc_buffer_0 vss vco_out vdd out_first_buffer out_to_div out_to_buffer ring_osc_buffer
Xdiv_by_5_0 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in n_out_by_2
+ div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/DFlipFlop_0/latch_diff_1/nD
+ vss vdd div_by_5_0/DFlipFlop_2/latch_diff_0/nD div_5_Q0 div_5_Q1 out_by_2 div_by_5_0/DFlipFlop_0/Q
+ div_by_5_0/DFlipFlop_2/latch_diff_1/D div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# div_5_nQ0 div_by_5_0/DFlipFlop_3/latch_diff_0/D
+ div_by_5_0/DFlipFlop_3/latch_diff_1/nD div_by_5_0/DFlipFlop_1/latch_diff_1/nD div_by_5_0/DFlipFlop_1/latch_diff_0/nD
+ div_by_5_0/DFlipFlop_1/latch_diff_0/D div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280#
+ out_div_by_5 div_5_Q1_shift div_5_nQ2 div_by_5_0/DFlipFlop_2/D div_by_5_0/DFlipFlop_2/latch_diff_1/nD
+ div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out div_by_5_0/DFlipFlop_1/latch_diff_1/D
+ div_by_5_0/DFlipFlop_1/D div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ div_by_5_0/DFlipFlop_0/latch_diff_0/nD div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368#
+ div_by_5_0/DFlipFlop_0/D div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_0/latch_diff_1/D div_by_5_0/DFlipFlop_2/nQ div_by_5_0/DFlipFlop_3/latch_diff_0/nD
+ div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out div_by_5_0/DFlipFlop_2/latch_diff_0/D
+ div_by_5_0/DFlipFlop_0/latch_diff_0/D div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ div_by_5_0/DFlipFlop_3/latch_diff_1/D div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368#
+ div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136#
+ div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_152_368# div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# div_by_5_0/DFlipFlop_3/nQ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136#
+ div_by_5
Xpfd_cp_interface_0 vss pfd_cp_interface_0/inverter_cp_x1_2/in vdd pfd_cp_interface_0/inverter_cp_x1_0/out
+ Down QA QB nDown Up nUp pfd_cp_interface
XPFD_0 vss vdd pfd_reset QB QA in_ref out_div_by_5 PFD
C0 vco_vctrl div_5_Q0 0.48fF
C1 n_out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/D 0.24fF
C2 out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/nD 0.23fF
C3 vco_vctrl vdd -1.02fF
C4 ring_osc_0/csvco_branch_2/cap_vco_0/t vdd 0.02fF
C5 vco_vctrl ring_osc_0/csvco_branch_2/vbp 0.26fF
C6 div_by_5_0/DFlipFlop_0/D vco_vctrl -0.45fF
C7 n_out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_1/nD 0.24fF
C8 div_5_nQ2 out_by_2 0.16fF
C9 out_to_div div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out -0.12fF
C10 out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.17fF
C11 n_out_by_2 div_5_Q1 1.04fF
C12 n_out_by_2 vco_vctrl 0.52fF
C13 out_by_2 div_5_Q0 0.09fF
C14 out_to_div vdd 0.21fF
C15 out_to_div div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in -0.16fF
C16 out_by_2 vdd 0.97fF
C17 vdd D0_vco 0.03fF
C18 n_out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/nD 0.24fF
C19 lf_vc vdd 0.02fF
C20 pswitch Up 1.98fF
C21 buffer_salida_0/a_678_n100# vdd 0.24fF
C22 div_by_5_0/DFlipFlop_0/latch_diff_1/D n_out_by_2 0.17fF
C23 div_by_5_0/DFlipFlop_0/D out_by_2 0.35fF
C24 nUp Up 2.72fF
C25 nUp vdd 0.05fF
C26 pfd_cp_interface_0/inverter_cp_x1_2/in vdd 0.01fF
C27 out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/D 0.23fF
C28 iref_cp vdd 0.15fF
C29 n_out_by_2 div_by_5_0/DFlipFlop_2/D 0.19fF
C30 n_out_by_2 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in -0.20fF
C31 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vdd 0.04fF
C32 nDown vdd 0.22fF
C33 biasp Up 0.26fF
C34 out_by_2 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out -0.04fF
C35 vco_vctrl div_5_Q1 0.14fF
C36 div_by_5_0/DFlipFlop_1/latch_diff_1/D out_by_2 0.23fF
C37 out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/D 0.09fF
C38 out_to_div out_to_buffer 0.13fF
C39 n_out_by_2 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.27fF
C40 n_out_by_2 div_by_5_0/DFlipFlop_0/Q -0.23fF
C41 out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_1/nD 0.09fF
C42 buffer_salida_0/a_678_n100# out_to_buffer 0.22fF
C43 n_out_by_2 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out -0.11fF
C44 vco_vctrl ring_osc_0/csvco_branch_0/inverter_csvco_0/vss 0.04fF
C45 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out out_by_2 0.28fF
C46 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# out_div_by_5 0.18fF
C47 out_by_2 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# 0.10fF
C48 out_div_by_5 vdd 0.28fF
C49 out_by_2 div_5_Q1 0.42fF
C50 n_out_by_2 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in -0.51fF
C51 div_5_Q1_shift out_div_by_5 0.05fF
C52 vco_vctrl out_by_2 0.53fF
C53 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# 0.03fF
C54 n_out_by_2 div_by_5_0/DFlipFlop_1/D 0.22fF
C55 out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/nD 0.09fF
C56 div_by_5_0/DFlipFlop_0/latch_diff_1/D out_by_2 0.33fF
C57 vco_vctrl nUp 0.02fF
C58 n_out_by_2 div_by_5_0/DFlipFlop_2/nQ 0.10fF
C59 n_out_by_2 div_5_nQ0 0.10fF
C60 out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_0/nD 0.10fF
C61 out_by_2 div_by_5_0/DFlipFlop_2/D 0.22fF
C62 n_out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_0/nD 0.11fF
C63 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# -0.05fF
C64 QA vdd -0.04fF
C65 out_by_2 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out 0.09fF
C66 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vdd 0.03fF
C67 out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_0/nD 0.10fF
C68 out_by_2 div_by_5_0/DFlipFlop_0/Q 0.09fF
C69 nswitch vco_vctrl -0.06fF
C70 n_out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/nD 0.10fF
C71 vdd Up 0.28fF
C72 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# 0.02fF
C73 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392# 0.01fF
C74 div_5_Q1 out_div_by_5 0.01fF
C75 pswitch nUp 0.85fF
C76 n_out_by_2 div_5_nQ2 0.10fF
C77 n_out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_0/D 0.12fF
C78 vdd ring_osc_0/csvco_branch_2/vbp 0.03fF
C79 pswitch nDown 0.53fF
C80 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# 0.12fF
C81 nUp nDown -0.09fF
C82 n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.33fF
C83 biasp nUp -0.17fF
C84 n_out_by_2 div_5_Q0 -0.12fF
C85 out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_0/D 0.11fF
C86 out_by_2 div_by_5_0/DFlipFlop_1/D 0.38fF
C87 iref_cp Down 0.09fF
C88 n_out_by_2 vdd 1.03fF
C89 biasp nDown 0.26fF
C90 n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_0/D 0.24fF
C91 nDown Down 2.55fF
C92 vco_vctrl div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# -0.11fF
C93 out_by_2 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in -0.22fF
C94 out_by_2 div_by_5_0/DFlipFlop_2/nQ 0.23fF
C95 div_5_nQ0 out_by_2 0.32fF
C96 biasp Down 1.24fF
C97 div_by_5_0/DFlipFlop_0/D n_out_by_2 -1.48fF
C98 vdd out_to_buffer 0.07fF
C99 n_out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_0/D 0.12fF
C100 out_first_buffer ring_osc_0/csvco_branch_2/cap_vco_0/t 0.03fF
C101 n_out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/D 0.10fF
C102 out_by_2 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136# -0.02fF
C103 nswitch nDown 0.76fF
C104 vco_vctrl div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# -0.36fF
C105 nswitch Down 0.54fF
C106 out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_0/nD 0.17fF
C107 n_out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_1/D 0.10fF
C108 PFD_0/and_pfd_0/a_656_410# vss 0.96fF
C109 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C110 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.07fF
C111 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C112 PFD_0/dff_pfd_1/nor_pfd_2/B vss 1.40fF
C113 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C114 PFD_0/dff_pfd_1/nor_pfd_3/A vss 3.14fF
C115 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C116 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C117 PFD_0/dff_pfd_1/nor_pfd_2/A vss 2.55fF
C118 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C119 QB vss 4.46fF
C120 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C121 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C122 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C123 out_div_by_5 vss -0.40fF
C124 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C125 PFD_0/dff_pfd_0/nor_pfd_2/B vss 1.40fF
C126 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C127 PFD_0/dff_pfd_0/nor_pfd_3/A vss 3.14fF
C128 pfd_reset vss 2.17fF
C129 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C130 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C131 PFD_0/dff_pfd_0/nor_pfd_2/A vss 2.55fF
C132 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C133 QA vss 4.31fF
C134 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C135 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C136 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C137 in_ref vss 1.19fF
C138 pfd_cp_interface_0/inverter_cp_x1_2/in vss 1.85fF
C139 pfd_cp_interface_0/inverter_cp_x1_0/out vss 1.87fF
C140 nUp vss 5.50fF
C141 Up vss 2.37fF
C142 Down vss 7.92fF
C143 nDown vss -2.20fF
C144 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C145 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.38fF
C146 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.41fF
C147 div_5_Q1_shift vss -0.14fF
C148 div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.57fF
C149 div_by_5_0/DFlipFlop_3/nQ vss 0.48fF
C150 div_by_5_0/DFlipFlop_3/latch_diff_1/D vss -1.73fF
C151 div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C152 div_by_5_0/DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C153 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C154 div_by_5_0/DFlipFlop_3/latch_diff_0/D vss 0.96fF
C155 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C156 div_by_5_0/DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C157 div_5_Q1 vss 4.28fF
C158 div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C159 div_by_5_0/DFlipFlop_2/nQ vss 0.48fF
C160 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C161 div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C162 div_by_5_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C163 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C164 div_by_5_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C165 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C166 div_by_5_0/DFlipFlop_2/D vss 3.13fF
C167 div_by_5_0/DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C168 div_5_Q0 vss 0.01fF
C169 div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C170 div_5_nQ0 vss 0.59fF
C171 div_by_5_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C172 div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C173 div_by_5_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C174 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C175 div_by_5_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C176 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C177 div_by_5_0/DFlipFlop_1/D vss 3.64fF
C178 div_by_5_0/DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C179 div_by_5_0/DFlipFlop_0/Q vss -0.94fF
C180 div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C181 n_out_by_2 vss -2.62fF
C182 div_5_nQ2 vss 1.24fF
C183 div_by_5_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C184 div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C185 out_by_2 vss -4.51fF
C186 div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C187 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C188 div_by_5_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C189 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C190 div_by_5_0/DFlipFlop_0/D vss 3.96fF
C191 vdd vss 366.82fF
C192 div_by_5_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C193 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C194 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.40fF
C195 out_first_buffer vss 2.88fF
C196 out_to_buffer vss 1.57fF
C197 out_to_div vss 4.46fF
C198 ring_osc_0/csvco_branch_2/in vss 1.60fF
C199 ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C200 ring_osc_0/csvco_branch_1/cap_vco_0/t vss 7.10fF
C201 ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vss 0.52fF
C202 ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C203 ring_osc_0/csvco_branch_2/cap_vco_0/t vss 7.10fF
C204 ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vss 0.52fF
C205 ring_osc_0/csvco_branch_1/in vss 1.58fF
C206 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C207 vco_out vss 1.01fF
C208 D0_vco vss -4.63fF
C209 ring_osc_0/csvco_branch_0/cap_vco_0/t vss 7.10fF
C210 ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vss 0.52fF
C211 ring_osc_0/csvco_branch_2/vbp vss 0.38fF
C212 out_to_pad vss 7.50fF
C213 buffer_salida_0/a_3996_n100# vss 48.29fF
C214 buffer_salida_0/a_678_n100# vss 13.38fF
C215 lf_vc vss -59.89fF
C216 loop_filter_v2_0/res_loop_filter_2/out vss 7.90fF
C217 DO_cap vss 0.01fF
C218 loop_filter_v2_0/cap3_loop_filter_0/in vss -12.03fF
C219 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C220 div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C221 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.89fF
C222 div_by_2_0/DFlipFlop_0/nCLK vss 1.03fF
C223 out_buffer_div_2 vss 1.60fF
C224 n_out_buffer_div_2 vss 1.63fF
C225 out_div_2 vss -1.30fF
C226 div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C227 div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C228 div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C229 div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C230 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C231 div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C232 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C233 n_out_div_2 vss 1.95fF
C234 div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C235 nswitch vss 3.73fF
C236 biasp vss 5.44fF
C237 iref_cp vss 2.81fF
C238 vco_vctrl vss -21.20fF
C239 pswitch vss 3.57fF
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xres_amp_top_0 vssa1 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_3/in
+ vdda1 bias_0/iref_9 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/a_3747_261# bias_0/iref_8
+ res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vp res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/out
+ bias_0/iref_6 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/in1
+ res_amp_top_0/res_amp_lin_prog_0/outn bias_0/iref_7 res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1384_n363#
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/out res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_pmos_0/m1_957_828#
+ gpio_noesd[3] bias_0/iref_5 res_amp_top_0/res_amp_lin_prog_0/outp res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/in
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/inverter_min_1/in
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinB io_analog[2]
+ res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_pmos_1/m1_957_828#
+ io_analog[3] res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_511_801# res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/sel_b
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_12/inverter_min_1/in
+ res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/clk res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinA
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/DinA gpio_noesd[1]
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_5/out res_amp_top_0/res_amp_lin_prog_0/outp_cap
+ gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/clk res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinB
+ res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/in res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vctrl
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_2/inverter_min_1/in
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinA io_analog[6]
+ gpio_noesd[5] res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_0/in
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/out gpio_noesd[6]
+ res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_964_n363# res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_10/inverter_min_1/in
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/out res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/sel_b
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/out res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/m1_21_n341#
+ res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_7/inverter_min_1/in
+ gpio_noesd[2] io_analog[0] res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/m1_460_n1129#
+ io_analog[1] io_analog[4] res_amp_top_0/res_amp_sync_v2_0/rst res_amp_top
Xtop_pll_v3_0 top_pll_v3_0/clk_d vdda1 gpio_noesd[10] top_pll_v3_0/charge_pump_0/w_2544_775#
+ top_pll_v3_0/out_by_2 top_pll_v3_0/s_0_n io_analog[10] top_pll_v3_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd
+ top_pll_v3_0/buffer_salida_0/a_3996_n100# vssa1 top_pll_v3_0/vco_vctrl gpio_noesd[9]
+ top_pll_v3_0/ring_osc_0/csvco_branch_2/vbp top_pll_v3_0/lf_vc gpio_noesd[7] gpio_noesd[8]
+ top_pll_v3_0/buffer_salida_0/a_678_n100# top_pll_v3_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd
+ top_pll_v3_0/loop_filter_v2_0/cap3_loop_filter_0/in top_pll_v3_0/charge_pump_0/w_1008_774#
+ bias_0/iref_0 top_pll_v3_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd top_pll_v3_0/Down
+ top_pll_v3_0/out_to_div top_pll_v3_0/clk_1 top_pll_v3_0/out_div top_pll_v3_0/nDown
+ top_pll_v3_0/s_1_n io_analog[7] gpio_noesd[11] top_pll_v3_0/Up top_pll_v3_0/clk_0
+ top_pll_v3_0/freq_div_0/prescaler_23_0/nCLK_23 top_pll_v3_0/biasp top_pll_v3_0/nUp
+ top_pll_v3_0/n_clk_0 top_pll_v3
Xtop_pll_v1_0 top_pll_v1_0/vco_vctrl top_pll_v1_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd
+ vdda1 top_pll_v1_0/charge_pump_0/w_2544_775# top_pll_v1_0/pswitch top_pll_v1_0/biasp
+ top_pll_v1_0/ring_osc_0/csvco_branch_2/vbp io_analog[10] top_pll_v1_0/Down vssa1
+ vssa1 gpio_noesd[7] top_pll_v1_0/QA top_pll_v1_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd
+ bias_0/iref_2 top_pll_v1_0/out_to_div top_pll_v1_0/nDown io_analog[9] top_pll_v1_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd
+ top_pll_v1_0/Up top_pll_v1_0/nUp top_pll_v1
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[0] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[1] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[2] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[3] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[4] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[5] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[6] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[7] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[8] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xbias_0 vssa1 vdda1 bias_0/iref_0 bias_0/iref_1 bias_0/iref_2 bias_0/iref_5 bias_0/iref_6
+ bias_0/iref_7 bias_0/iref_8 bias_0/iref_9 io_analog[5] bias
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[0] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[1] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[2] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[3] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[4] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[5] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[6] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[7] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[8] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xmimcap_decoup_1x5_0[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_0[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_0[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_1[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_1[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_1[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[0] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[1] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[2] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[3] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[4] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[5] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[6] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xmimcap_decoup_1x5_2[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_2[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_2[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_3[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_3[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_3[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_4[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_4[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_4[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_5[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_5[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_5[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_6[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_6[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xtop_pll_v2_0 top_pll_v2_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd top_pll_v2_0/pswitch
+ vdda1 top_pll_v2_0/charge_pump_0/w_2544_775# top_pll_v2_0/ring_osc_0/csvco_branch_2/vbp
+ top_pll_v2_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd io_analog[10] top_pll_v2_0/vco_vctrl
+ top_pll_v2_0/Down vssa1 vssa1 gpio_noesd[7] bias_0/iref_1 top_pll_v2_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd
+ top_pll_v2_0/out_to_div gpio_noesd[8] top_pll_v2_0/nDown top_pll_v2_0/biasp io_analog[8]
+ top_pll_v2_0/Up top_pll_v2_0/nUp top_pll_v2
C0 vdda1 gpio_noesd[9] 65.72fF
C1 top_pll_v3_0/clk_1 gpio_noesd[10] 0.49fF
C2 vdda1 top_pll_v2_0/pswitch 0.34fF
C3 gpio_noesd[1] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_2/inverter_min_1/in 0.18fF
C4 vdda1 top_pll_v2_0/ring_osc_0/csvco_branch_2/vbp 2.10fF
C5 gpio_noesd[4] io_analog[3] -0.78fF
C6 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_pmos_1/m1_957_828# bias_0/iref_8 0.11fF
C7 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/m1_460_n1129# bias_0/iref_6 0.15fF
C8 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/DinA gpio_noesd[1] 0.29fF
C9 bias_0/iref_2 io_analog[8] 14.44fF
C10 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinA gpio_noesd[2] 0.72fF
C11 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/inverter_min_1/in gpio_noesd[5] 0.05fF
C12 io_analog[2] gpio_noesd[5] 0.09fF
C13 vdda1 top_pll_v2_0/nUp 0.01fF
C14 vdda1 io_analog[0] 76.77fF
C15 bias_0/iref_1 top_pll_v2_0/nDown 0.54fF
C16 vdda1 io_analog[9] 30.05fF
C17 bias_0/iref_2 top_pll_v1_0/nDown 0.70fF
C18 top_pll_v3_0/lf_vc gpio_noesd[10] 0.48fF
C19 gpio_noesd[4] bias_0/iref_9 -0.25fF
C20 io_analog[4] bias_0/iref_6 15.97fF
C21 res_amp_top_0/res_amp_lin_prog_0/outn gpio_noesd[5] 1.42fF
C22 bias_0/iref_2 top_pll_v1_0/charge_pump_0/w_2544_775# 0.02fF
C23 vdda1 top_pll_v2_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd 0.17fF
C24 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/out gpio_noesd[2] 0.21fF
C25 io_analog[10] top_pll_v1_0/QA 0.03fF
C26 vdda1 top_pll_v1_0/ring_osc_0/csvco_branch_2/vbp 1.01fF
C27 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_5/out gpio_noesd[3] 0.33fF
C28 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/clk gpio_noesd[6] 2.12fF
C29 gpio_noesd[9] gpio_noesd[11] 0.96fF
C30 top_pll_v3_0/out_to_div gpio_noesd[7] 4.28fF
C31 gpio_noesd[6] res_amp_top_0/res_amp_lin_prog_0/outp 0.61fF
C32 vdda1 top_pll_v3_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd 0.12fF
C33 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/m1_460_n1129# bias_0/iref_5 0.45fF
C34 bias_0/iref_2 io_analog[9] 14.44fF
C35 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/in gpio_noesd[5] 0.47fF
C36 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinA gpio_noesd[3] 0.01fF
C37 gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_964_n363# -0.11fF
C38 vdda1 top_pll_v1_0/nUp 0.01fF
C39 bias_0/iref_9 res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1384_n363# 0.78fF
C40 gpio_noesd[1] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/out 0.57fF
C41 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vp gpio_noesd[5] 0.54fF
C42 vdda1 top_pll_v1_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd 0.04fF
C43 bias_0/iref_1 top_pll_v2_0/Up 0.54fF
C44 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/out gpio_noesd[3] 0.03fF
C45 io_analog[4] bias_0/iref_5 15.97fF
C46 gpio_noesd[1] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/out 0.21fF
C47 vdda1 io_analog[3] 25.90fF
C48 bias_0/iref_2 top_pll_v1_0/nUp 0.70fF
C49 gpio_noesd[10] top_pll_v3_0/out_by_2 0.10fF
C50 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vctrl gpio_noesd[5] 0.33fF
C51 gpio_noesd[7] top_pll_v2_0/vco_vctrl 0.05fF
C52 vdda1 top_pll_v2_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd 0.17fF
C53 vdda1 bias_0/iref_7 33.08fF
C54 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/a_3747_261# gpio_noesd[5] 0.14fF
C55 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinB gpio_noesd[5] 0.14fF
C56 vdda1 bias_0/iref_9 30.24fF
C57 io_analog[10] gpio_noesd[7] 29.88fF
C58 io_analog[6] io_clamp_high[2] 0.53fF
C59 top_pll_v1_0/vco_vctrl gpio_noesd[7] 0.05fF
C60 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/out gpio_noesd[2] 0.38fF
C61 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/clk gpio_noesd[4] -0.13fF
C62 bias_0/iref_1 top_pll_v2_0/biasp 2.20fF
C63 vdda1 gpio_noesd[6] 53.94fF
C64 gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/outp -0.31fF
C65 bias_0/iref_5 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/in 0.46fF
C66 top_pll_v3_0/vco_vctrl gpio_noesd[10] 0.53fF
C67 io_analog[4] io_clamp_high[0] 0.53fF
C68 vdda1 top_pll_v1_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd 0.04fF
C69 res_amp_top_0/res_amp_lin_prog_0/clk gpio_noesd[4] -0.01fF
C70 io_clamp_low[2] io_clamp_high[2] 0.53fF
C71 vdda1 bias_0/iref_8 31.37fF
C72 top_pll_v3_0/lf_vc gpio_noesd[8] 2.98fF
C73 io_analog[3] bias_0/iref_6 13.88fF
C74 gpio_noesd[3] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_10/inverter_min_1/in -0.70fF
C75 bias_0/iref_0 top_pll_v3_0/charge_pump_0/w_2544_775# 0.21fF
C76 vdda1 top_pll_v2_0/biasp 0.03fF
C77 bias_0/iref_7 bias_0/iref_6 17.40fF
C78 bias_0/iref_7 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_0/in 0.94fF
C79 bias_0/iref_0 top_pll_v3_0/Up 0.74fF
C80 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/m1_21_n341# gpio_noesd[5] 0.16fF
C81 gpio_noesd[9] io_analog[10] 1.87fF
C82 vdda1 gpio_noesd[10] 53.94fF
C83 vdda1 gpio_noesd[4] 117.64fF
C84 gpio_noesd[3] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinB 0.01fF
C85 io_analog[3] bias_0/iref_5 13.88fF
C86 bias_0/iref_1 top_pll_v2_0/Down 0.91fF
C87 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/in1 gpio_noesd[5] 0.26fF
C88 io_analog[2] io_analog[3] 0.14fF
C89 io_clamp_low[1] io_clamp_high[1] 0.53fF
C90 bias_0/iref_7 bias_0/iref_5 10.35fF
C91 io_analog[2] bias_0/iref_7 13.88fF
C92 bias_0/iref_0 top_pll_v3_0/nUp 0.74fF
C93 io_analog[6] gpio_noesd[10] 25.05fF
C94 vdda1 bias_0/iref_1 15.26fF
C95 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/out gpio_noesd[2] 0.21fF
C96 io_analog[2] bias_0/iref_9 13.88fF
C97 vdda1 top_pll_v1_0/biasp 0.03fF
C98 io_analog[3] gpio_noesd[5] 0.12fF
C99 gpio_noesd[10] top_pll_v3_0/freq_div_0/prescaler_23_0/nCLK_23 1.35fF
C100 vdda1 top_pll_v3_0/buffer_salida_0/a_3996_n100# 1.78fF
C101 io_analog[5] io_clamp_high[1] 0.53fF
C102 gpio_noesd[1] res_amp_top_0/res_amp_lin_prog_0/clk 0.39fF
C103 gpio_noesd[10] gpio_noesd[11] 39.51fF
C104 bias_0/iref_8 bias_0/iref_5 10.19fF
C105 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_5/out gpio_noesd[4] 0.19fF
C106 io_analog[2] bias_0/iref_8 13.88fF
C107 io_analog[6] bias_0/iref_1 13.22fF
C108 bias_0/iref_2 top_pll_v1_0/biasp 3.20fF
C109 bias_0/iref_9 gpio_noesd[5] 1.30fF
C110 gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_12/inverter_min_1/in 0.12fF
C111 gpio_noesd[6] res_amp_top_0/res_amp_lin_prog_0/outn 0.45fF
C112 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinA gpio_noesd[4] 0.42fF
C113 io_analog[7] bias_0/iref_1 13.22fF
C114 gpio_noesd[6] gpio_noesd[5] 0.05fF
C115 top_pll_v3_0/buffer_salida_0/a_3996_n100# io_analog[7] -0.08fF
C116 gpio_noesd[10] top_pll_v3_0/s_0_n 0.31fF
C117 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinB gpio_noesd[2] 0.19fF
C118 bias_0/iref_7 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/m1_460_n1129# 0.45fF
C119 vdda1 top_pll_v2_0/buffer_salida_0/a_3996_n100# 0.05fF
C120 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_pmos_0/m1_957_828# bias_0/iref_7 0.09fF
C121 vdda1 top_pll_v3_0/buffer_salida_0/a_678_n100# 0.50fF
C122 vdda1 bias_0/iref_2 3.90fF
C123 bias_0/iref_9 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vctrl 0.42fF
C124 vdda1 top_pll_v3_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd 0.12fF
C125 vdda1 io_analog[6] 124.15fF
C126 vdda1 gpio_noesd[8] 77.43fF
C127 gpio_noesd[10] top_pll_v3_0/clk_0 0.12fF
C128 bias_0/iref_2 top_pll_v1_0/Down 1.11fF
C129 vdda1 gpio_noesd[1] 214.54fF
C130 io_analog[4] bias_0/iref_7 15.97fF
C131 vdda1 io_analog[7] 29.48fF
C132 gpio_noesd[6] res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vctrl 0.22fF
C133 gpio_noesd[9] top_pll_v3_0/clk_d 0.15fF
C134 io_clamp_low[0] io_clamp_high[0] 0.53fF
C135 gpio_noesd[4] io_analog[2] -0.21fF
C136 vdda1 gpio_noesd[11] 102.31fF
C137 vdda1 top_pll_v1_0/pswitch 0.38fF
C138 vdda1 top_pll_v1_0/buffer_salida_0/a_3996_n100# 0.06fF
C139 io_analog[4] bias_0/iref_9 15.97fF
C140 io_analog[6] bias_0/iref_2 54.67fF
C141 vdda1 top_pll_v3_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd 0.12fF
C142 bias_0/iref_0 top_pll_v3_0/nDown 0.74fF
C143 io_analog[7] bias_0/iref_2 13.22fF
C144 gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/outn -1.06fF
C145 vdda1 bias_0/iref_6 29.75fF
C146 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/clk gpio_noesd[5] 0.44fF
C147 gpio_noesd[4] gpio_noesd[5] 4.67fF
C148 bias_0/iref_2 top_pll_v1_0/Up 0.70fF
C149 res_amp_top_0/res_amp_lin_prog_0/outp gpio_noesd[5] 0.44fF
C150 io_analog[4] bias_0/iref_8 15.97fF
C151 io_analog[6] gpio_noesd[11] 9.16fF
C152 bias_0/iref_7 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/in 1.46fF
C153 io_analog[6] io_clamp_low[2] 0.53fF
C154 res_amp_top_0/res_amp_lin_prog_0/clk gpio_noesd[5] 0.68fF
C155 gpio_noesd[11] top_pll_v3_0/freq_div_0/prescaler_23_0/nCLK_23 0.17fF
C156 vdda1 top_pll_v2_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd 0.17fF
C157 gpio_noesd[2] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinA 0.49fF
C158 gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vp 0.17fF
C159 io_analog[4] io_clamp_low[0] 0.53fF
C160 top_pll_v3_0/vco_vctrl gpio_noesd[7] 0.13fF
C161 gpio_noesd[5] res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1384_n363# 0.32fF
C162 res_amp_top_0/res_amp_lin_prog_0/outp_cap bias_0/iref_7 0.37fF
C163 gpio_noesd[1] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_3/in 0.23fF
C164 gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vctrl 0.07fF
C165 gpio_noesd[10] io_analog[10] 1.87fF
C166 vdda1 bias_0/iref_5 30.67fF
C167 bias_0/iref_8 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/in 1.34fF
C168 vdda1 io_analog[2] 25.90fF
C169 gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/a_3747_261# -0.08fF
C170 vdda1 top_pll_v1_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd 0.04fF
C171 res_amp_top_0/res_amp_lin_prog_0/clk gpio_noesd[2] 0.37fF
C172 gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinB 0.08fF
C173 top_pll_v3_0/loop_filter_v2_0/cap3_loop_filter_0/in gpio_noesd[8] 3.13fF
C174 vdda1 io_analog[1] 76.56fF
C175 res_amp_top_0/res_amp_lin_prog_0/outp_cap bias_0/iref_8 0.37fF
C176 bias_0/iref_0 top_pll_v3_0/Down 1.08fF
C177 vdda1 gpio_noesd[5] 124.75fF
C178 bias_0/iref_1 top_pll_v2_0/charge_pump_0/w_2544_775# 0.09fF
C179 gpio_noesd[2] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/sel_b 0.31fF
C180 io_analog[3] bias_0/iref_7 13.88fF
C181 vdda1 top_pll_v3_0/ring_osc_0/csvco_branch_2/vbp 1.07fF
C182 vdda1 gpio_noesd[7] 120.96fF
C183 gpio_noesd[10] gpio_noesd[9] 0.96fF
C184 bias_0/iref_0 top_pll_v3_0/charge_pump_0/w_1008_774# 0.21fF
C185 vdda1 top_pll_v2_0/vco_vctrl 0.59fF
C186 io_analog[3] bias_0/iref_9 13.88fF
C187 res_amp_top_0/res_amp_lin_prog_0/clk gpio_noesd[3] 0.21fF
C188 bias_0/iref_0 vdda1 15.18fF
C189 gpio_noesd[10] top_pll_v3_0/n_clk_0 0.10fF
C190 bias_0/iref_5 bias_0/iref_6 29.11fF
C191 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_0/in bias_0/iref_5 0.46fF
C192 gpio_noesd[7] top_pll_v2_0/out_to_div 0.23fF
C193 vdda1 io_analog[10] 0.01fF
C194 io_analog[2] bias_0/iref_6 13.88fF
C195 vdda1 top_pll_v1_0/vco_vctrl 0.43fF
C196 gpio_noesd[4] res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_511_801# 0.18fF
C197 io_analog[3] bias_0/iref_8 13.88fF
C198 gpio_noesd[8] gpio_noesd[7] 5.92fF
C199 vdda1 gpio_noesd[2] 214.16fF
C200 bias_0/iref_7 bias_0/iref_8 13.23fF
C201 bias_0/iref_0 io_analog[6] 6.93fF
C202 io_analog[5] io_clamp_low[1] 0.53fF
C203 gpio_noesd[2] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_7/inverter_min_1/in 0.20fF
C204 vdda1 io_analog[4] 182.26fF
C205 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_pmos_1/m1_957_828# bias_0/iref_7 0.40fF
C206 gpio_noesd[9] top_pll_v3_0/out_div 0.16fF
C207 top_pll_v3_0/s_1_n gpio_noesd[9] 0.08fF
C208 gpio_noesd[8] io_analog[10] 20.65fF
C209 bias_0/iref_9 bias_0/iref_8 9.89fF
C210 bias_0/iref_0 top_pll_v3_0/biasp 3.13fF
C211 gpio_noesd[1] res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/sel_b 0.23fF
C212 top_pll_v1_0/out_to_div gpio_noesd[7] 0.23fF
C213 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/in1 gpio_noesd[4] -0.05fF
C214 bias_0/iref_1 top_pll_v2_0/nUp 0.22fF
C215 res_amp_top_0/res_amp_sync_v2_0/rst bias_0/iref_9 0.39fF
C216 gpio_noesd[1] gpio_noesd[2] 0.30fF
C217 bias_0/iref_5 io_analog[5] 0.09fF
C218 io_analog[2] bias_0/iref_5 13.88fF
C219 vdda1 gpio_noesd[3] 120.88fF
C220 gpio_noesd[11] io_analog[10] 1.87fF
C221 vdda1 io_analog[8] 29.93fF
C222 io_analog[6] io_analog[4] 0.59fF
C223 io_in_3v3[0] vssa1 0.41fF
C224 io_oeb[26] vssa1 0.61fF
C225 io_in[0] vssa1 0.41fF
C226 io_out[26] vssa1 0.61fF
C227 io_out[0] vssa1 0.41fF
C228 io_in[26] vssa1 0.61fF
C229 io_oeb[0] vssa1 0.41fF
C230 io_in_3v3[26] vssa1 0.61fF
C231 io_in_3v3[1] vssa1 0.41fF
C232 io_oeb[25] vssa1 0.61fF
C233 io_in[1] vssa1 0.41fF
C234 io_out[25] vssa1 0.61fF
C235 io_out[1] vssa1 0.41fF
C236 io_in[25] vssa1 0.61fF
C237 io_oeb[1] vssa1 0.41fF
C238 io_in_3v3[25] vssa1 0.61fF
C239 io_in_3v3[2] vssa1 0.41fF
C240 io_oeb[24] vssa1 0.61fF
C241 io_in[2] vssa1 0.41fF
C242 io_out[24] vssa1 0.61fF
C243 io_out[2] vssa1 0.41fF
C244 io_in[24] vssa1 0.61fF
C245 io_oeb[2] vssa1 -0.20fF
C246 io_in_3v3[3] vssa1 0.41fF
C247 gpio_noesd[17] vssa1 0.61fF
C248 io_in[3] vssa1 0.41fF
C249 gpio_analog[17] vssa1 0.61fF
C250 io_out[3] vssa1 0.41fF
C251 io_oeb[3] vssa1 0.41fF
C252 io_in_3v3[4] vssa1 0.41fF
C253 io_in[4] vssa1 0.41fF
C254 io_out[4] vssa1 0.41fF
C255 io_oeb[4] vssa1 0.41fF
C256 io_oeb[23] vssa1 0.61fF
C257 io_out[23] vssa1 0.61fF
C258 io_in[23] vssa1 0.61fF
C259 io_in_3v3[23] vssa1 0.61fF
C260 gpio_noesd[16] vssa1 0.61fF
C261 io_in_3v3[5] vssa1 0.41fF
C262 io_in[5] vssa1 -0.20fF
C263 io_out[5] vssa1 0.41fF
C264 io_oeb[5] vssa1 0.41fF
C265 io_oeb[22] vssa1 0.61fF
C266 io_out[22] vssa1 0.61fF
C267 io_in[22] vssa1 0.61fF
C268 io_in_3v3[22] vssa1 0.61fF
C269 gpio_analog[15] vssa1 0.61fF
C270 io_in_3v3[6] vssa1 -0.20fF
C271 io_in[6] vssa1 0.41fF
C272 io_out[6] vssa1 0.41fF
C273 io_oeb[6] vssa1 0.41fF
C274 io_oeb[21] vssa1 0.61fF
C275 io_out[21] vssa1 0.61fF
C276 io_in[21] vssa1 0.61fF
C277 io_in_3v3[21] vssa1 0.61fF
C278 gpio_noesd[14] vssa1 0.61fF
C279 gpio_analog[14] vssa1 0.61fF
C280 vssd2 vssa1 -5.19fF
C281 vssd1 vssa1 1.13fF
C282 vdda2 vssa1 -5.19fF
C283 io_oeb[20] vssa1 0.61fF
C284 io_out[20] vssa1 0.61fF
C285 io_in[20] vssa1 0.61fF
C286 io_in_3v3[20] vssa1 0.61fF
C287 gpio_noesd[13] vssa1 0.61fF
C288 gpio_analog[13] vssa1 0.61fF
C289 gpio_analog[0] vssa1 0.41fF
C290 gpio_noesd[0] vssa1 0.41fF
C291 io_in_3v3[7] vssa1 0.41fF
C292 io_in[7] vssa1 0.41fF
C293 io_out[7] vssa1 0.41fF
C294 io_oeb[7] vssa1 0.41fF
C295 io_oeb[19] vssa1 0.61fF
C296 io_out[19] vssa1 0.61fF
C297 io_in[19] vssa1 0.61fF
C298 io_in_3v3[19] vssa1 0.61fF
C299 gpio_noesd[12] vssa1 0.61fF
C300 gpio_analog[12] vssa1 0.61fF
C301 gpio_analog[1] vssa1 0.41fF
C302 io_in_3v3[8] vssa1 0.41fF
C303 io_in[8] vssa1 0.41fF
C304 io_out[8] vssa1 -0.20fF
C305 io_oeb[8] vssa1 0.41fF
C306 gpio_analog[2] vssa1 0.41fF
C307 io_in_3v3[9] vssa1 0.41fF
C308 io_in[9] vssa1 0.41fF
C309 io_out[9] vssa1 0.41fF
C310 io_oeb[9] vssa1 0.41fF
C311 gpio_analog[3] vssa1 0.41fF
C312 io_in_3v3[10] vssa1 0.41fF
C313 io_in[10] vssa1 0.41fF
C314 io_out[10] vssa1 0.41fF
C315 io_oeb[10] vssa1 0.41fF
C316 gpio_analog[4] vssa1 0.41fF
C317 io_in_3v3[11] vssa1 0.41fF
C318 io_in[11] vssa1 0.41fF
C319 io_out[11] vssa1 0.41fF
C320 io_oeb[11] vssa1 0.41fF
C321 gpio_analog[5] vssa1 0.41fF
C322 io_in_3v3[12] vssa1 0.41fF
C323 io_in[12] vssa1 0.41fF
C324 io_out[12] vssa1 0.41fF
C325 io_oeb[12] vssa1 0.41fF
C326 gpio_analog[6] vssa1 0.60fF
C327 io_in_3v3[13] vssa1 0.60fF
C328 io_in[13] vssa1 0.60fF
C329 io_out[13] vssa1 0.60fF
C330 io_oeb[13] vssa1 0.60fF
C331 io_oeb[18] vssa1 0.61fF
C332 io_out[18] vssa1 0.61fF
C333 io_in_3v3[18] vssa1 0.61fF
C334 vccd1 vssa1 0.85fF
C335 gpio_analog[11] vssa1 0.61fF
C336 io_oeb[17] vssa1 0.61fF
C337 io_in[17] vssa1 0.61fF
C338 io_in_3v3[17] vssa1 0.61fF
C339 gpio_analog[10] vssa1 0.61fF
C340 io_out[16] vssa1 0.61fF
C341 io_in[16] vssa1 0.61fF
C342 io_in_3v3[16] vssa1 0.61fF
C343 gpio_analog[9] vssa1 0.61fF
C344 io_oeb[15] vssa1 0.61fF
C345 io_out[15] vssa1 0.61fF
C346 io_in[15] vssa1 0.61fF
C347 io_in_3v3[15] vssa1 0.61fF
C348 gpio_analog[8] vssa1 0.61fF
C349 io_oeb[14] vssa1 0.61fF
C350 io_out[14] vssa1 0.61fF
C351 io_in[14] vssa1 0.61fF
C352 io_in_3v3[14] vssa1 0.61fF
C353 vssa2 vssa1 1.66fF
C354 vccd2 vssa1 0.91fF
C355 io_clamp_high[0] vssa1 -2.60fF
C356 io_clamp_low[0] vssa1 0.82fF
C357 io_clamp_high[1] vssa1 0.71fF
C358 io_clamp_low[1] vssa1 0.55fF
C359 io_clamp_high[2] vssa1 0.66fF
C360 io_clamp_low[2] vssa1 0.50fF
C361 user_irq[2] vssa1 0.63fF
C362 user_irq[1] vssa1 0.63fF
C363 user_irq[0] vssa1 0.63fF
C364 user_clock2 vssa1 0.63fF
C365 la_oenb[127] vssa1 0.63fF
C366 la_data_in[127] vssa1 0.63fF
C367 la_oenb[126] vssa1 0.63fF
C368 la_data_out[126] vssa1 0.63fF
C369 la_data_in[126] vssa1 0.63fF
C370 la_oenb[125] vssa1 0.63fF
C371 la_data_out[125] vssa1 0.63fF
C372 la_data_in[125] vssa1 0.63fF
C373 la_oenb[124] vssa1 0.63fF
C374 la_data_out[124] vssa1 0.63fF
C375 la_data_in[124] vssa1 0.63fF
C376 la_oenb[123] vssa1 0.63fF
C377 la_data_out[123] vssa1 0.63fF
C378 la_oenb[122] vssa1 0.63fF
C379 la_data_out[122] vssa1 0.63fF
C380 la_data_in[122] vssa1 0.63fF
C381 la_oenb[121] vssa1 0.63fF
C382 la_data_out[121] vssa1 0.63fF
C383 la_data_in[121] vssa1 0.63fF
C384 la_oenb[120] vssa1 0.63fF
C385 la_data_out[120] vssa1 0.63fF
C386 la_data_in[120] vssa1 0.63fF
C387 la_oenb[119] vssa1 0.63fF
C388 la_data_out[119] vssa1 0.63fF
C389 la_data_in[119] vssa1 0.63fF
C390 la_oenb[118] vssa1 0.63fF
C391 la_data_out[118] vssa1 0.63fF
C392 la_data_in[118] vssa1 0.63fF
C393 la_oenb[117] vssa1 0.63fF
C394 la_data_out[117] vssa1 0.63fF
C395 la_data_in[117] vssa1 0.63fF
C396 la_data_out[116] vssa1 0.63fF
C397 la_data_in[116] vssa1 0.63fF
C398 la_oenb[115] vssa1 0.63fF
C399 la_data_out[115] vssa1 0.63fF
C400 la_data_in[115] vssa1 0.63fF
C401 la_oenb[114] vssa1 0.63fF
C402 la_data_out[114] vssa1 0.63fF
C403 la_data_in[114] vssa1 0.63fF
C404 la_oenb[113] vssa1 0.63fF
C405 la_data_out[113] vssa1 0.63fF
C406 la_data_in[113] vssa1 0.63fF
C407 la_oenb[112] vssa1 0.63fF
C408 la_data_in[112] vssa1 0.63fF
C409 la_oenb[111] vssa1 0.63fF
C410 la_data_out[111] vssa1 0.63fF
C411 la_data_in[111] vssa1 0.63fF
C412 la_oenb[110] vssa1 0.63fF
C413 la_data_out[110] vssa1 0.63fF
C414 la_data_in[110] vssa1 0.63fF
C415 la_oenb[109] vssa1 0.63fF
C416 la_data_out[109] vssa1 0.63fF
C417 la_data_in[109] vssa1 0.63fF
C418 la_oenb[108] vssa1 0.63fF
C419 la_data_out[108] vssa1 0.63fF
C420 la_oenb[107] vssa1 0.63fF
C421 la_data_out[107] vssa1 0.63fF
C422 la_data_in[107] vssa1 0.63fF
C423 la_oenb[106] vssa1 0.63fF
C424 la_data_out[106] vssa1 0.63fF
C425 la_oenb[105] vssa1 0.63fF
C426 la_data_out[105] vssa1 0.63fF
C427 la_data_in[105] vssa1 0.63fF
C428 la_oenb[104] vssa1 0.63fF
C429 la_data_out[104] vssa1 0.63fF
C430 la_data_in[104] vssa1 0.63fF
C431 la_oenb[103] vssa1 0.63fF
C432 la_data_out[103] vssa1 0.63fF
C433 la_data_in[103] vssa1 0.63fF
C434 la_oenb[102] vssa1 0.63fF
C435 la_data_out[102] vssa1 0.63fF
C436 la_data_in[102] vssa1 0.63fF
C437 la_data_out[101] vssa1 0.63fF
C438 la_data_in[101] vssa1 0.63fF
C439 la_oenb[100] vssa1 0.63fF
C440 la_data_out[100] vssa1 0.63fF
C441 la_data_in[100] vssa1 0.63fF
C442 la_oenb[99] vssa1 0.63fF
C443 la_data_out[99] vssa1 0.63fF
C444 la_data_in[99] vssa1 0.63fF
C445 la_oenb[98] vssa1 0.63fF
C446 la_data_out[98] vssa1 0.63fF
C447 la_data_in[98] vssa1 0.63fF
C448 la_oenb[97] vssa1 0.63fF
C449 la_data_in[97] vssa1 0.63fF
C450 la_oenb[96] vssa1 0.63fF
C451 la_data_out[96] vssa1 0.63fF
C452 la_data_in[96] vssa1 0.63fF
C453 la_oenb[95] vssa1 0.63fF
C454 la_data_out[95] vssa1 0.63fF
C455 la_data_in[95] vssa1 0.63fF
C456 la_oenb[94] vssa1 0.63fF
C457 la_data_out[94] vssa1 0.63fF
C458 la_data_in[94] vssa1 0.63fF
C459 la_oenb[93] vssa1 0.63fF
C460 la_data_out[93] vssa1 0.63fF
C461 la_oenb[92] vssa1 0.63fF
C462 la_data_out[92] vssa1 0.63fF
C463 la_data_in[92] vssa1 0.63fF
C464 la_oenb[91] vssa1 0.63fF
C465 la_data_out[91] vssa1 0.63fF
C466 la_oenb[90] vssa1 0.63fF
C467 la_data_out[90] vssa1 0.63fF
C468 la_data_in[90] vssa1 0.63fF
C469 la_oenb[89] vssa1 0.63fF
C470 la_data_out[89] vssa1 0.63fF
C471 la_data_in[89] vssa1 0.63fF
C472 la_oenb[88] vssa1 0.63fF
C473 la_data_out[88] vssa1 0.63fF
C474 la_data_in[88] vssa1 0.63fF
C475 la_oenb[87] vssa1 0.63fF
C476 la_data_out[87] vssa1 0.63fF
C477 la_data_in[87] vssa1 0.63fF
C478 la_data_out[86] vssa1 0.63fF
C479 la_data_in[86] vssa1 0.63fF
C480 la_oenb[85] vssa1 0.63fF
C481 la_data_out[85] vssa1 0.63fF
C482 la_data_in[85] vssa1 0.63fF
C483 la_oenb[84] vssa1 0.63fF
C484 la_data_out[84] vssa1 0.63fF
C485 la_data_in[84] vssa1 0.63fF
C486 la_oenb[83] vssa1 0.63fF
C487 la_data_out[83] vssa1 0.63fF
C488 la_data_in[83] vssa1 0.63fF
C489 la_oenb[82] vssa1 0.63fF
C490 la_data_in[82] vssa1 0.63fF
C491 la_oenb[81] vssa1 0.63fF
C492 la_data_out[81] vssa1 0.63fF
C493 la_data_in[81] vssa1 0.63fF
C494 la_oenb[80] vssa1 0.63fF
C495 la_data_out[80] vssa1 0.63fF
C496 la_data_in[80] vssa1 0.63fF
C497 la_oenb[79] vssa1 0.63fF
C498 la_data_out[79] vssa1 0.63fF
C499 la_data_in[79] vssa1 0.63fF
C500 la_oenb[78] vssa1 0.63fF
C501 la_data_out[78] vssa1 0.63fF
C502 la_data_in[78] vssa1 0.63fF
C503 la_oenb[77] vssa1 0.63fF
C504 la_data_out[77] vssa1 0.63fF
C505 la_data_in[77] vssa1 0.63fF
C506 la_oenb[76] vssa1 0.63fF
C507 la_data_out[76] vssa1 0.63fF
C508 la_oenb[75] vssa1 0.63fF
C509 la_data_out[75] vssa1 0.63fF
C510 la_data_in[75] vssa1 0.63fF
C511 la_oenb[74] vssa1 0.63fF
C512 la_data_out[74] vssa1 0.63fF
C513 la_data_in[74] vssa1 0.63fF
C514 la_oenb[73] vssa1 0.63fF
C515 la_data_out[73] vssa1 0.63fF
C516 la_data_in[73] vssa1 0.63fF
C517 la_oenb[72] vssa1 0.63fF
C518 la_data_out[72] vssa1 0.63fF
C519 la_data_in[72] vssa1 0.63fF
C520 la_data_out[71] vssa1 0.63fF
C521 la_data_in[71] vssa1 0.63fF
C522 la_oenb[70] vssa1 0.63fF
C523 la_data_out[70] vssa1 0.63fF
C524 la_data_in[70] vssa1 0.63fF
C525 la_oenb[69] vssa1 0.63fF
C526 la_data_out[69] vssa1 0.63fF
C527 la_data_in[69] vssa1 0.63fF
C528 la_oenb[68] vssa1 0.63fF
C529 la_data_out[68] vssa1 0.63fF
C530 la_data_in[68] vssa1 0.63fF
C531 la_oenb[67] vssa1 0.63fF
C532 la_data_in[67] vssa1 0.63fF
C533 la_oenb[66] vssa1 0.63fF
C534 la_data_out[66] vssa1 0.63fF
C535 la_data_in[66] vssa1 0.63fF
C536 la_oenb[65] vssa1 0.63fF
C537 la_data_out[65] vssa1 0.26fF
C538 la_data_in[65] vssa1 0.63fF
C539 la_oenb[64] vssa1 0.63fF
C540 la_data_out[64] vssa1 0.63fF
C541 la_data_in[64] vssa1 0.63fF
C542 la_oenb[63] vssa1 0.63fF
C543 la_data_out[63] vssa1 0.63fF
C544 la_data_in[63] vssa1 0.63fF
C545 la_oenb[62] vssa1 0.63fF
C546 la_data_out[62] vssa1 0.63fF
C547 la_data_in[62] vssa1 0.63fF
C548 la_oenb[61] vssa1 0.63fF
C549 la_data_out[61] vssa1 0.63fF
C550 la_oenb[60] vssa1 0.63fF
C551 la_data_out[60] vssa1 0.63fF
C552 la_data_in[60] vssa1 0.63fF
C553 la_oenb[59] vssa1 0.63fF
C554 la_data_out[59] vssa1 0.63fF
C555 la_data_in[59] vssa1 0.63fF
C556 la_oenb[58] vssa1 0.63fF
C557 la_data_out[58] vssa1 0.63fF
C558 la_data_in[58] vssa1 0.63fF
C559 la_oenb[57] vssa1 0.63fF
C560 la_data_out[57] vssa1 0.63fF
C561 la_data_in[57] vssa1 0.63fF
C562 la_data_out[56] vssa1 0.63fF
C563 la_data_in[56] vssa1 0.63fF
C564 la_oenb[55] vssa1 0.63fF
C565 la_data_out[55] vssa1 0.63fF
C566 la_data_in[55] vssa1 0.63fF
C567 la_oenb[54] vssa1 0.63fF
C568 la_data_out[54] vssa1 0.63fF
C569 la_data_in[54] vssa1 0.63fF
C570 la_oenb[53] vssa1 0.63fF
C571 la_data_out[53] vssa1 0.63fF
C572 la_data_in[53] vssa1 0.63fF
C573 la_oenb[52] vssa1 0.63fF
C574 la_data_in[52] vssa1 0.63fF
C575 la_oenb[51] vssa1 0.63fF
C576 la_data_out[51] vssa1 0.63fF
C577 la_data_in[51] vssa1 0.63fF
C578 la_oenb[50] vssa1 0.63fF
C579 la_data_in[50] vssa1 0.63fF
C580 la_oenb[49] vssa1 0.63fF
C581 la_data_out[49] vssa1 0.63fF
C582 la_data_in[49] vssa1 0.63fF
C583 la_oenb[48] vssa1 0.63fF
C584 la_data_out[48] vssa1 0.63fF
C585 la_data_in[48] vssa1 0.63fF
C586 la_oenb[47] vssa1 0.63fF
C587 la_data_out[47] vssa1 0.63fF
C588 la_data_in[47] vssa1 0.63fF
C589 la_oenb[46] vssa1 0.63fF
C590 la_data_out[46] vssa1 0.63fF
C591 la_oenb[45] vssa1 0.63fF
C592 la_data_out[45] vssa1 0.63fF
C593 la_data_in[45] vssa1 0.63fF
C594 la_oenb[44] vssa1 0.63fF
C595 la_data_out[44] vssa1 0.63fF
C596 la_data_in[44] vssa1 0.63fF
C597 la_oenb[43] vssa1 0.63fF
C598 la_data_out[43] vssa1 0.63fF
C599 la_data_in[43] vssa1 0.63fF
C600 la_oenb[42] vssa1 0.63fF
C601 la_data_out[42] vssa1 0.63fF
C602 la_data_in[42] vssa1 0.63fF
C603 la_data_out[41] vssa1 0.63fF
C604 la_data_in[41] vssa1 0.63fF
C605 la_oenb[40] vssa1 0.63fF
C606 la_data_out[40] vssa1 0.63fF
C607 la_data_in[40] vssa1 0.63fF
C608 la_oenb[39] vssa1 0.63fF
C609 la_data_out[39] vssa1 0.63fF
C610 la_data_in[39] vssa1 0.63fF
C611 la_oenb[38] vssa1 0.63fF
C612 la_data_out[38] vssa1 0.63fF
C613 la_data_in[38] vssa1 0.63fF
C614 la_oenb[37] vssa1 0.63fF
C615 la_data_out[37] vssa1 0.26fF
C616 la_data_in[37] vssa1 0.63fF
C617 la_oenb[36] vssa1 0.63fF
C618 la_data_out[36] vssa1 0.63fF
C619 la_data_in[36] vssa1 0.63fF
C620 la_oenb[35] vssa1 0.63fF
C621 la_data_in[35] vssa1 0.63fF
C622 la_oenb[34] vssa1 0.63fF
C623 la_data_out[34] vssa1 0.63fF
C624 la_data_in[34] vssa1 0.63fF
C625 la_oenb[33] vssa1 0.63fF
C626 la_data_out[33] vssa1 0.63fF
C627 la_data_in[33] vssa1 0.63fF
C628 la_oenb[32] vssa1 0.63fF
C629 la_data_out[32] vssa1 0.63fF
C630 la_data_in[32] vssa1 0.63fF
C631 la_oenb[31] vssa1 0.63fF
C632 la_data_out[31] vssa1 0.63fF
C633 la_oenb[30] vssa1 0.63fF
C634 la_data_out[30] vssa1 0.63fF
C635 la_data_in[30] vssa1 0.63fF
C636 la_oenb[29] vssa1 0.63fF
C637 la_data_out[29] vssa1 0.63fF
C638 la_data_in[29] vssa1 0.63fF
C639 la_oenb[28] vssa1 0.63fF
C640 la_data_out[28] vssa1 0.63fF
C641 la_data_in[28] vssa1 0.63fF
C642 la_oenb[27] vssa1 0.63fF
C643 la_data_out[27] vssa1 0.63fF
C644 la_data_in[27] vssa1 0.63fF
C645 la_data_out[26] vssa1 0.63fF
C646 la_data_in[26] vssa1 0.63fF
C647 la_oenb[25] vssa1 0.63fF
C648 la_data_out[25] vssa1 0.63fF
C649 la_data_in[25] vssa1 0.63fF
C650 la_oenb[24] vssa1 0.63fF
C651 la_data_out[24] vssa1 0.63fF
C652 la_data_in[24] vssa1 0.63fF
C653 la_oenb[23] vssa1 0.63fF
C654 la_data_out[23] vssa1 0.63fF
C655 la_data_in[23] vssa1 0.63fF
C656 la_oenb[22] vssa1 0.63fF
C657 la_data_out[22] vssa1 0.63fF
C658 la_data_in[22] vssa1 0.63fF
C659 la_oenb[21] vssa1 0.63fF
C660 la_data_out[21] vssa1 0.63fF
C661 la_data_in[21] vssa1 0.63fF
C662 la_oenb[20] vssa1 0.63fF
C663 la_data_in[20] vssa1 0.63fF
C664 la_oenb[19] vssa1 0.63fF
C665 la_data_out[19] vssa1 0.63fF
C666 la_data_in[19] vssa1 0.63fF
C667 la_oenb[18] vssa1 0.63fF
C668 la_data_out[18] vssa1 0.63fF
C669 la_data_in[18] vssa1 0.63fF
C670 la_oenb[17] vssa1 0.63fF
C671 la_data_out[17] vssa1 0.63fF
C672 la_data_in[17] vssa1 0.63fF
C673 la_oenb[16] vssa1 0.63fF
C674 la_data_out[16] vssa1 0.63fF
C675 la_oenb[15] vssa1 0.63fF
C676 la_data_out[15] vssa1 0.63fF
C677 la_data_in[15] vssa1 0.63fF
C678 la_oenb[14] vssa1 0.63fF
C679 la_data_out[14] vssa1 0.63fF
C680 la_data_in[14] vssa1 0.63fF
C681 la_oenb[13] vssa1 0.63fF
C682 la_data_out[13] vssa1 0.63fF
C683 la_data_in[13] vssa1 0.63fF
C684 la_oenb[12] vssa1 0.63fF
C685 la_data_out[12] vssa1 0.63fF
C686 la_data_in[12] vssa1 0.63fF
C687 la_data_out[11] vssa1 0.63fF
C688 la_data_in[11] vssa1 0.63fF
C689 la_oenb[10] vssa1 0.63fF
C690 la_data_out[10] vssa1 0.63fF
C691 la_data_in[10] vssa1 0.63fF
C692 la_data_out[9] vssa1 0.63fF
C693 la_data_in[9] vssa1 0.63fF
C694 la_oenb[8] vssa1 0.63fF
C695 la_data_out[8] vssa1 0.63fF
C696 la_data_in[8] vssa1 0.63fF
C697 la_oenb[7] vssa1 0.63fF
C698 la_data_out[7] vssa1 0.63fF
C699 la_data_in[7] vssa1 0.63fF
C700 la_oenb[6] vssa1 0.63fF
C701 la_data_out[6] vssa1 0.63fF
C702 la_data_in[6] vssa1 0.63fF
C703 la_oenb[5] vssa1 0.63fF
C704 la_data_in[5] vssa1 0.63fF
C705 la_oenb[4] vssa1 0.63fF
C706 la_data_out[4] vssa1 0.63fF
C707 la_data_in[4] vssa1 0.63fF
C708 la_oenb[3] vssa1 0.63fF
C709 la_data_out[3] vssa1 0.63fF
C710 la_data_in[3] vssa1 0.63fF
C711 la_oenb[2] vssa1 0.63fF
C712 la_data_out[2] vssa1 0.63fF
C713 la_data_in[2] vssa1 0.63fF
C714 la_oenb[1] vssa1 0.63fF
C715 la_data_out[1] vssa1 0.63fF
C716 la_oenb[0] vssa1 0.63fF
C717 la_data_out[0] vssa1 0.63fF
C718 la_data_in[0] vssa1 0.63fF
C719 wbs_dat_o[31] vssa1 0.63fF
C720 wbs_dat_i[31] vssa1 0.63fF
C721 wbs_adr_i[31] vssa1 0.63fF
C722 wbs_dat_o[30] vssa1 0.63fF
C723 wbs_dat_i[30] vssa1 0.63fF
C724 wbs_adr_i[30] vssa1 0.63fF
C725 wbs_dat_o[29] vssa1 0.63fF
C726 wbs_dat_i[29] vssa1 0.63fF
C727 wbs_adr_i[29] vssa1 0.63fF
C728 wbs_dat_i[28] vssa1 0.63fF
C729 wbs_adr_i[28] vssa1 0.63fF
C730 wbs_dat_o[27] vssa1 0.63fF
C731 wbs_dat_i[27] vssa1 0.63fF
C732 wbs_adr_i[27] vssa1 0.63fF
C733 wbs_dat_i[26] vssa1 0.63fF
C734 wbs_adr_i[26] vssa1 0.63fF
C735 wbs_dat_o[25] vssa1 0.63fF
C736 wbs_dat_i[25] vssa1 0.63fF
C737 wbs_adr_i[25] vssa1 0.63fF
C738 wbs_dat_o[24] vssa1 0.63fF
C739 wbs_dat_i[24] vssa1 0.63fF
C740 wbs_adr_i[24] vssa1 0.63fF
C741 wbs_dat_o[23] vssa1 0.63fF
C742 wbs_dat_i[23] vssa1 0.63fF
C743 wbs_adr_i[23] vssa1 0.63fF
C744 wbs_dat_o[22] vssa1 0.63fF
C745 wbs_adr_i[22] vssa1 0.63fF
C746 wbs_dat_o[21] vssa1 0.63fF
C747 wbs_dat_i[21] vssa1 0.63fF
C748 wbs_adr_i[21] vssa1 0.63fF
C749 wbs_dat_o[20] vssa1 0.63fF
C750 wbs_dat_i[20] vssa1 0.63fF
C751 wbs_adr_i[20] vssa1 0.63fF
C752 wbs_dat_o[19] vssa1 0.63fF
C753 wbs_dat_i[19] vssa1 0.63fF
C754 wbs_adr_i[19] vssa1 0.63fF
C755 wbs_dat_o[18] vssa1 0.63fF
C756 wbs_dat_i[18] vssa1 0.63fF
C757 wbs_dat_o[17] vssa1 0.63fF
C758 wbs_dat_i[17] vssa1 0.63fF
C759 wbs_adr_i[17] vssa1 0.63fF
C760 wbs_dat_o[16] vssa1 0.63fF
C761 wbs_dat_i[16] vssa1 0.63fF
C762 wbs_adr_i[16] vssa1 0.63fF
C763 wbs_dat_o[15] vssa1 0.63fF
C764 wbs_dat_i[15] vssa1 0.63fF
C765 wbs_adr_i[15] vssa1 0.63fF
C766 wbs_dat_o[14] vssa1 0.63fF
C767 wbs_dat_i[14] vssa1 0.63fF
C768 wbs_adr_i[14] vssa1 0.63fF
C769 wbs_dat_o[13] vssa1 0.63fF
C770 wbs_dat_i[13] vssa1 0.63fF
C771 wbs_adr_i[13] vssa1 0.63fF
C772 wbs_dat_o[12] vssa1 0.63fF
C773 wbs_dat_i[12] vssa1 0.63fF
C774 wbs_adr_i[12] vssa1 0.63fF
C775 wbs_dat_i[11] vssa1 0.63fF
C776 wbs_adr_i[11] vssa1 0.63fF
C777 wbs_dat_o[10] vssa1 0.63fF
C778 wbs_dat_i[10] vssa1 0.63fF
C779 wbs_adr_i[10] vssa1 0.63fF
C780 wbs_dat_o[9] vssa1 0.63fF
C781 wbs_dat_i[9] vssa1 0.63fF
C782 wbs_adr_i[9] vssa1 0.63fF
C783 wbs_dat_o[8] vssa1 0.63fF
C784 wbs_dat_i[8] vssa1 0.63fF
C785 wbs_adr_i[8] vssa1 0.63fF
C786 wbs_dat_o[7] vssa1 0.63fF
C787 wbs_adr_i[7] vssa1 0.63fF
C788 wbs_dat_o[6] vssa1 0.63fF
C789 wbs_dat_i[6] vssa1 0.63fF
C790 wbs_adr_i[6] vssa1 0.63fF
C791 wbs_dat_o[5] vssa1 0.63fF
C792 wbs_dat_i[5] vssa1 0.63fF
C793 wbs_adr_i[5] vssa1 0.63fF
C794 wbs_dat_o[4] vssa1 0.63fF
C795 wbs_dat_i[4] vssa1 0.63fF
C796 wbs_adr_i[4] vssa1 0.63fF
C797 wbs_sel_i[3] vssa1 0.63fF
C798 wbs_dat_o[3] vssa1 0.63fF
C799 wbs_adr_i[3] vssa1 0.63fF
C800 wbs_sel_i[2] vssa1 0.63fF
C801 wbs_dat_o[2] vssa1 0.63fF
C802 wbs_dat_i[2] vssa1 0.63fF
C803 wbs_adr_i[2] vssa1 0.63fF
C804 wbs_dat_o[1] vssa1 0.63fF
C805 wbs_dat_i[1] vssa1 0.63fF
C806 wbs_adr_i[1] vssa1 0.63fF
C807 wbs_sel_i[0] vssa1 0.63fF
C808 wbs_dat_o[0] vssa1 0.63fF
C809 wbs_dat_i[0] vssa1 0.63fF
C810 wbs_adr_i[0] vssa1 0.63fF
C811 wbs_we_i vssa1 0.63fF
C812 wbs_stb_i vssa1 0.63fF
C813 wbs_cyc_i vssa1 0.63fF
C814 wbs_ack_o vssa1 0.63fF
C815 wb_rst_i vssa1 0.63fF
C816 top_pll_v2_0/PFD_0/and_pfd_0/a_656_410# vssa1 0.96fF
C817 top_pll_v2_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vssa1 0.05fF
C818 top_pll_v2_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vssa1 0.05fF
C819 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C820 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_2/B vssa1 1.40fF
C821 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C822 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_3/A vssa1 3.14fF
C823 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C824 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C825 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_2/A vssa1 2.55fF
C826 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C827 top_pll_v2_0/QB vssa1 4.35fF
C828 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C829 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C830 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C831 top_pll_v2_0/out_div_by_5 vssa1 -0.40fF
C832 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C833 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_2/B vssa1 1.40fF
C834 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C835 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_3/A vssa1 3.14fF
C836 top_pll_v2_0/pfd_reset vssa1 2.17fF
C837 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C838 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C839 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_2/A vssa1 2.55fF
C840 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C841 top_pll_v2_0/QA vssa1 4.22fF
C842 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C843 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C844 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C845 top_pll_v2_0/pfd_cp_interface_0/inverter_cp_x1_2/in vssa1 1.85fF
C846 top_pll_v2_0/pfd_cp_interface_0/inverter_cp_x1_0/out vssa1 1.77fF
C847 top_pll_v2_0/nUp vssa1 5.39fF
C848 top_pll_v2_0/Up vssa1 1.85fF
C849 top_pll_v2_0/Down vssa1 6.19fF
C850 top_pll_v2_0/nDown vssa1 -3.53fF
C851 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vssa1 0.37fF
C852 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vssa1 0.38fF
C853 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vssa1 0.38fF
C854 top_pll_v2_0/div_5_Q1_shift vssa1 -0.14fF
C855 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vssa1 0.57fF
C856 top_pll_v2_0/div_by_5_0/DFlipFlop_3/nQ vssa1 0.48fF
C857 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_1/D vssa1 -1.73fF
C858 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vssa1 0.57fF
C859 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_1/nD vssa1 0.57fF
C860 top_pll_v2_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C861 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_0/D vssa1 0.96fF
C862 top_pll_v2_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C863 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_0/nD vssa1 1.14fF
C864 top_pll_v2_0/div_5_Q1 vssa1 4.25fF
C865 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vssa1 0.57fF
C866 top_pll_v2_0/div_by_5_0/DFlipFlop_2/nQ vssa1 0.48fF
C867 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D vssa1 -1.73fF
C868 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vssa1 0.57fF
C869 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD vssa1 0.57fF
C870 top_pll_v2_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C871 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D vssa1 0.96fF
C872 top_pll_v2_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C873 top_pll_v2_0/div_by_5_0/DFlipFlop_2/D vssa1 3.13fF
C874 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD vssa1 1.14fF
C875 top_pll_v2_0/div_5_Q0 vssa1 0.01fF
C876 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vssa1 0.57fF
C877 top_pll_v2_0/div_5_nQ0 vssa1 0.59fF
C878 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_1/D vssa1 -1.73fF
C879 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vssa1 0.57fF
C880 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_1/nD vssa1 0.57fF
C881 top_pll_v2_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C882 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_0/D vssa1 0.96fF
C883 top_pll_v2_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C884 top_pll_v2_0/div_by_5_0/DFlipFlop_1/D vssa1 3.64fF
C885 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_0/nD vssa1 1.14fF
C886 top_pll_v2_0/div_by_5_0/DFlipFlop_0/Q vssa1 -0.94fF
C887 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C888 top_pll_v2_0/n_out_by_2 vssa1 -2.75fF
C889 top_pll_v2_0/div_5_nQ2 vssa1 1.24fF
C890 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C891 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C892 top_pll_v2_0/out_by_2 vssa1 -5.01fF
C893 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C894 top_pll_v2_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C895 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C896 top_pll_v2_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C897 top_pll_v2_0/div_by_5_0/DFlipFlop_0/D vssa1 3.96fF
C898 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C899 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vssa1 0.08fF
C900 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vssa1 0.40fF
C901 top_pll_v2_0/out_first_buffer vssa1 2.88fF
C902 top_pll_v2_0/out_to_buffer vssa1 1.54fF
C903 top_pll_v2_0/out_to_div vssa1 4.23fF
C904 top_pll_v2_0/ring_osc_0/csvco_branch_2/in vssa1 1.60fF
C905 top_pll_v2_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vssa1 0.16fF
C906 top_pll_v2_0/ring_osc_0/csvco_branch_1/cap_vco_0/t vssa1 7.10fF
C907 top_pll_v2_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vssa1 0.52fF
C908 top_pll_v2_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vssa1 0.16fF
C909 top_pll_v2_0/ring_osc_0/csvco_branch_2/cap_vco_0/t vssa1 7.10fF
C910 top_pll_v2_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vssa1 0.52fF
C911 top_pll_v2_0/ring_osc_0/csvco_branch_1/in vssa1 1.58fF
C912 top_pll_v2_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vssa1 0.16fF
C913 top_pll_v2_0/vco_out vssa1 1.01fF
C914 top_pll_v2_0/ring_osc_0/csvco_branch_0/cap_vco_0/t vssa1 7.10fF
C915 top_pll_v2_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vssa1 0.52fF
C916 top_pll_v2_0/ring_osc_0/csvco_branch_2/vbp vssa1 0.36fF
C917 io_analog[8] vssa1 13.78fF
C918 top_pll_v2_0/buffer_salida_0/a_3996_n100# vssa1 48.23fF
C919 top_pll_v2_0/buffer_salida_0/a_678_n100# vssa1 13.21fF
C920 top_pll_v2_0/lf_vc vssa1 -59.89fF
C921 top_pll_v2_0/loop_filter_v2_0/res_loop_filter_2/out vssa1 7.90fF
C922 top_pll_v2_0/loop_filter_v2_0/cap3_loop_filter_0/in vssa1 -12.03fF
C923 top_pll_v2_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C924 top_pll_v2_0/div_by_2_0/DFlipFlop_0/CLK vssa1 0.31fF
C925 top_pll_v2_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C926 top_pll_v2_0/div_by_2_0/DFlipFlop_0/nCLK vssa1 1.03fF
C927 top_pll_v2_0/out_buffer_div_2 vssa1 1.60fF
C928 top_pll_v2_0/n_out_buffer_div_2 vssa1 1.63fF
C929 top_pll_v2_0/out_div_2 vssa1 -1.30fF
C930 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C931 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C932 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C933 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C934 top_pll_v2_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C935 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C936 top_pll_v2_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C937 top_pll_v2_0/n_out_div_2 vssa1 1.95fF
C938 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C939 top_pll_v2_0/nswitch vssa1 3.73fF
C940 top_pll_v2_0/biasp vssa1 5.44fF
C941 bias_0/iref_1 vssa1 -91.53fF
C942 top_pll_v2_0/vco_vctrl vssa1 -20.08fF
C943 top_pll_v2_0/pswitch vssa1 3.57fF
C944 bias_0/iref_4 vssa1 1.17fF
C945 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# vssa1 2.60fF
C946 bias_0/iref_3 vssa1 0.64fF
C947 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# vssa1 2.60fF
C948 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219# vssa1 2.60fF
C949 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# vssa1 2.60fF
C950 io_analog[5] vssa1 33.29fF
C951 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_0/a_n1731_n1219# vssa1 2.60fF
C952 bias_0/m1_20168_984# vssa1 56.92fF
C953 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219# vssa1 2.60fF
C954 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219# vssa1 2.60fF
C955 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219# vssa1 2.60fF
C956 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219# vssa1 2.60fF
C957 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_6/a_n1731_n1219# vssa1 2.60fF
C958 top_pll_v1_0/PFD_0/and_pfd_0/a_656_410# vssa1 0.96fF
C959 top_pll_v1_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vssa1 0.05fF
C960 top_pll_v1_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vssa1 0.05fF
C961 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C962 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_2/B vssa1 1.40fF
C963 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C964 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_3/A vssa1 3.14fF
C965 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C966 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C967 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_2/A vssa1 2.55fF
C968 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C969 top_pll_v1_0/QB vssa1 4.35fF
C970 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C971 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C972 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C973 top_pll_v1_0/out_div_by_5 vssa1 -0.40fF
C974 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C975 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_2/B vssa1 1.40fF
C976 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C977 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_3/A vssa1 3.14fF
C978 top_pll_v1_0/pfd_reset vssa1 2.17fF
C979 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C980 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C981 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_2/A vssa1 2.55fF
C982 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C983 top_pll_v1_0/QA vssa1 4.22fF
C984 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C985 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C986 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C987 top_pll_v1_0/pfd_cp_interface_0/inverter_cp_x1_2/in vssa1 1.85fF
C988 top_pll_v1_0/pfd_cp_interface_0/inverter_cp_x1_0/out vssa1 1.77fF
C989 top_pll_v1_0/nUp vssa1 5.39fF
C990 top_pll_v1_0/Up vssa1 1.85fF
C991 top_pll_v1_0/Down vssa1 6.19fF
C992 top_pll_v1_0/nDown vssa1 -3.53fF
C993 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vssa1 0.37fF
C994 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vssa1 0.38fF
C995 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vssa1 0.38fF
C996 top_pll_v1_0/div_5_Q1_shift vssa1 -0.14fF
C997 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vssa1 0.57fF
C998 top_pll_v1_0/div_by_5_0/DFlipFlop_3/nQ vssa1 0.48fF
C999 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_1/D vssa1 -1.73fF
C1000 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vssa1 0.57fF
C1001 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_1/nD vssa1 0.57fF
C1002 top_pll_v1_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1003 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_0/D vssa1 0.96fF
C1004 top_pll_v1_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1005 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_0/nD vssa1 1.14fF
C1006 top_pll_v1_0/div_5_Q1 vssa1 4.25fF
C1007 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vssa1 0.57fF
C1008 top_pll_v1_0/div_by_5_0/DFlipFlop_2/nQ vssa1 0.48fF
C1009 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D vssa1 -1.73fF
C1010 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vssa1 0.57fF
C1011 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD vssa1 0.57fF
C1012 top_pll_v1_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1013 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D vssa1 0.96fF
C1014 top_pll_v1_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1015 top_pll_v1_0/div_by_5_0/DFlipFlop_2/D vssa1 3.13fF
C1016 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD vssa1 1.14fF
C1017 top_pll_v1_0/div_5_Q0 vssa1 0.01fF
C1018 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vssa1 0.57fF
C1019 top_pll_v1_0/div_5_nQ0 vssa1 0.59fF
C1020 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_1/D vssa1 -1.73fF
C1021 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vssa1 0.57fF
C1022 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_1/nD vssa1 0.57fF
C1023 top_pll_v1_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1024 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_0/D vssa1 0.96fF
C1025 top_pll_v1_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1026 top_pll_v1_0/div_by_5_0/DFlipFlop_1/D vssa1 3.64fF
C1027 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_0/nD vssa1 1.14fF
C1028 top_pll_v1_0/div_by_5_0/DFlipFlop_0/Q vssa1 -0.94fF
C1029 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C1030 top_pll_v1_0/n_out_by_2 vssa1 -2.75fF
C1031 top_pll_v1_0/div_5_nQ2 vssa1 1.24fF
C1032 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C1033 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C1034 top_pll_v1_0/out_by_2 vssa1 -5.01fF
C1035 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C1036 top_pll_v1_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1037 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C1038 top_pll_v1_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1039 top_pll_v1_0/div_by_5_0/DFlipFlop_0/D vssa1 3.96fF
C1040 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C1041 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vssa1 0.08fF
C1042 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vssa1 0.40fF
C1043 top_pll_v1_0/out_first_buffer vssa1 2.88fF
C1044 top_pll_v1_0/out_to_buffer vssa1 1.54fF
C1045 top_pll_v1_0/out_to_div vssa1 4.23fF
C1046 top_pll_v1_0/ring_osc_0/csvco_branch_2/in vssa1 1.60fF
C1047 top_pll_v1_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vssa1 0.16fF
C1048 top_pll_v1_0/ring_osc_0/csvco_branch_1/cap_vco_0/t vssa1 7.10fF
C1049 top_pll_v1_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vssa1 0.52fF
C1050 top_pll_v1_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vssa1 0.16fF
C1051 top_pll_v1_0/ring_osc_0/csvco_branch_2/cap_vco_0/t vssa1 7.10fF
C1052 top_pll_v1_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vssa1 0.52fF
C1053 top_pll_v1_0/ring_osc_0/csvco_branch_1/in vssa1 1.58fF
C1054 top_pll_v1_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vssa1 0.16fF
C1055 top_pll_v1_0/vco_out vssa1 1.01fF
C1056 gpio_noesd[7] vssa1 271.92fF
C1057 top_pll_v1_0/ring_osc_0/csvco_branch_0/cap_vco_0/t vssa1 7.10fF
C1058 top_pll_v1_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vssa1 0.52fF
C1059 top_pll_v1_0/ring_osc_0/csvco_branch_2/vbp vssa1 0.36fF
C1060 io_analog[9] vssa1 7.89fF
C1061 top_pll_v1_0/buffer_salida_0/a_3996_n100# vssa1 48.23fF
C1062 top_pll_v1_0/buffer_salida_0/a_678_n100# vssa1 13.21fF
C1063 top_pll_v1_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1064 top_pll_v1_0/div_by_2_0/DFlipFlop_0/CLK vssa1 0.31fF
C1065 top_pll_v1_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1066 top_pll_v1_0/div_by_2_0/DFlipFlop_0/nCLK vssa1 1.03fF
C1067 top_pll_v1_0/out_buffer_div_2 vssa1 1.60fF
C1068 top_pll_v1_0/n_out_buffer_div_2 vssa1 1.63fF
C1069 top_pll_v1_0/out_div_2 vssa1 -1.30fF
C1070 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C1071 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C1072 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C1073 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C1074 top_pll_v1_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1075 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C1076 top_pll_v1_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1077 top_pll_v1_0/n_out_div_2 vssa1 1.95fF
C1078 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C1079 top_pll_v1_0/nswitch vssa1 3.73fF
C1080 top_pll_v1_0/biasp vssa1 5.44fF
C1081 bias_0/iref_2 vssa1 -178.91fF
C1082 top_pll_v1_0/vco_vctrl vssa1 -18.17fF
C1083 top_pll_v1_0/pswitch vssa1 3.57fF
C1084 top_pll_v1_0/lf_vc vssa1 -59.89fF
C1085 top_pll_v1_0/loop_filter_0/res_loop_filter_2/out vssa1 7.90fF
C1086 top_pll_v3_0/PFD_0/and_pfd_0/a_656_410# vssa1 0.96fF
C1087 top_pll_v3_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vssa1 0.05fF
C1088 top_pll_v3_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vssa1 0.05fF
C1089 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C1090 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_2/B vssa1 1.40fF
C1091 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C1092 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_3/A vssa1 3.14fF
C1093 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C1094 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C1095 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_2/A vssa1 2.55fF
C1096 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C1097 top_pll_v3_0/QB vssa1 3.01fF
C1098 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C1099 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C1100 top_pll_v3_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C1101 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C1102 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_2/B vssa1 1.40fF
C1103 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C1104 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_3/A vssa1 3.14fF
C1105 top_pll_v3_0/pfd_reset vssa1 1.87fF
C1106 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C1107 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C1108 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_2/A vssa1 2.55fF
C1109 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C1110 top_pll_v3_0/QA vssa1 3.41fF
C1111 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C1112 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C1113 top_pll_v3_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C1114 io_analog[10] vssa1 502.98fF
C1115 top_pll_v3_0/pfd_cp_interface_0/inverter_cp_x1_2/in vssa1 1.85fF
C1116 top_pll_v3_0/pfd_cp_interface_0/inverter_cp_x1_0/out vssa1 1.77fF
C1117 top_pll_v3_0/Up vssa1 -4.79fF
C1118 top_pll_v3_0/Down vssa1 -0.05fF
C1119 top_pll_v3_0/nDown vssa1 1.54fF
C1120 top_pll_v3_0/out_first_buffer vssa1 2.14fF
C1121 top_pll_v3_0/out_to_buffer vssa1 1.89fF
C1122 top_pll_v3_0/out_to_div vssa1 8.23fF
C1123 top_pll_v3_0/ring_osc_0/csvco_branch_2/in vssa1 1.60fF
C1124 top_pll_v3_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vssa1 0.16fF
C1125 top_pll_v3_0/ring_osc_0/csvco_branch_1/cap_vco_0/t vssa1 7.10fF
C1126 top_pll_v3_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vssa1 0.52fF
C1127 top_pll_v3_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vssa1 0.16fF
C1128 top_pll_v3_0/ring_osc_0/csvco_branch_2/cap_vco_0/t vssa1 7.10fF
C1129 top_pll_v3_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vssa1 0.52fF
C1130 top_pll_v3_0/ring_osc_0/csvco_branch_1/in vssa1 1.58fF
C1131 top_pll_v3_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vssa1 0.16fF
C1132 top_pll_v3_0/vco_out vssa1 1.65fF
C1133 top_pll_v3_0/ring_osc_0/csvco_branch_0/cap_vco_0/t vssa1 7.10fF
C1134 top_pll_v3_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vssa1 0.52fF
C1135 top_pll_v3_0/ring_osc_0/csvco_branch_2/vbp vssa1 0.36fF
C1136 top_pll_v3_0/freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_1/a_63_368# vssa1 0.37fF
C1137 top_pll_v3_0/freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vssa1 0.37fF
C1138 top_pll_v3_0/freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_0/X vssa1 0.49fF
C1139 top_pll_v3_0/freq_div_0/prescaler_23_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vssa1 0.38fF
C1140 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_1/m1_657_280# vssa1 0.57fF
C1141 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_1/D vssa1 -1.73fF
C1142 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_0/m1_657_280# vssa1 0.57fF
C1143 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_1/nD vssa1 0.57fF
C1144 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1145 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_0/D vssa1 0.96fF
C1146 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1147 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_1/D vssa1 1.90fF
C1148 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_0/nD vssa1 1.14fF
C1149 top_pll_v3_0/freq_div_0/prescaler_23_0/Q2_d vssa1 -0.69fF
C1150 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# vssa1 0.57fF
C1151 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_2/nQ vssa1 0.48fF
C1152 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/D vssa1 -1.73fF
C1153 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# vssa1 0.57fF
C1154 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/nD vssa1 0.57fF
C1155 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1156 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/D vssa1 0.96fF
C1157 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1158 top_pll_v3_0/freq_div_0/prescaler_23_0/Q2 vssa1 0.55fF
C1159 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/nD vssa1 1.14fF
C1160 top_pll_v3_0/freq_div_0/prescaler_23_0/Q1 vssa1 0.07fF
C1161 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C1162 top_pll_v3_0/n_clk_0 vssa1 -7.01fF
C1163 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_0/nQ vssa1 0.48fF
C1164 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C1165 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C1166 top_pll_v3_0/clk_0 vssa1 -0.37fF
C1167 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C1168 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1169 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C1170 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1171 top_pll_v3_0/freq_div_0/prescaler_23_0/nCLK_23 vssa1 -1.02fF
C1172 top_pll_v3_0/freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C1173 top_pll_v3_0/freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_1/X vssa1 -1.01fF
C1174 gpio_noesd[11] vssa1 104.40fF
C1175 top_pll_v3_0/freq_div_0/prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_304_74# vssa1 0.36fF
C1176 top_pll_v3_0/freq_div_0/prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_27_112# vssa1 0.65fF
C1177 top_pll_v3_0/n_out_by_2 vssa1 4.38fF
C1178 top_pll_v3_0/s_0_n vssa1 -4.09fF
C1179 top_pll_v3_0/out_by_2 vssa1 4.28fF
C1180 gpio_noesd[10] vssa1 110.89fF
C1181 top_pll_v3_0/freq_div_0/div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vssa1 0.37fF
C1182 top_pll_v3_0/freq_div_0/div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vssa1 0.38fF
C1183 top_pll_v3_0/freq_div_0/div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vssa1 0.38fF
C1184 top_pll_v3_0/freq_div_0/div_by_5_0/Q1_shift vssa1 -0.36fF
C1185 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vssa1 0.57fF
C1186 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_3/nQ vssa1 0.48fF
C1187 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_1/D vssa1 -1.73fF
C1188 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vssa1 0.57fF
C1189 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_1/nD vssa1 0.57fF
C1190 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1191 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_0/D vssa1 0.96fF
C1192 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1193 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_0/nD vssa1 1.14fF
C1194 top_pll_v3_0/freq_div_0/div_by_5_0/Q1 vssa1 4.35fF
C1195 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vssa1 0.57fF
C1196 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/nQ vssa1 0.48fF
C1197 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D vssa1 -1.73fF
C1198 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vssa1 0.57fF
C1199 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD vssa1 0.57fF
C1200 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1201 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D vssa1 0.96fF
C1202 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1203 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/D vssa1 3.13fF
C1204 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD vssa1 1.14fF
C1205 top_pll_v3_0/freq_div_0/div_by_5_0/Q0 vssa1 0.29fF
C1206 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vssa1 0.57fF
C1207 top_pll_v3_0/freq_div_0/div_by_5_0/nQ0 vssa1 0.99fF
C1208 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_1/D vssa1 -1.73fF
C1209 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vssa1 0.57fF
C1210 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_1/nD vssa1 0.57fF
C1211 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1212 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_0/D vssa1 0.96fF
C1213 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1214 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_1/D vssa1 3.64fF
C1215 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_0/nD vssa1 1.14fF
C1216 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/Q vssa1 -0.94fF
C1217 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C1218 top_pll_v3_0/n_clk_1 vssa1 -0.56fF
C1219 top_pll_v3_0/freq_div_0/div_by_5_0/nQ2 vssa1 1.38fF
C1220 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C1221 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C1222 top_pll_v3_0/clk_1 vssa1 -2.08fF
C1223 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C1224 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1225 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C1226 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1227 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/D vssa1 3.96fF
C1228 top_pll_v3_0/freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C1229 top_pll_v3_0/freq_div_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vssa1 0.08fF
C1230 top_pll_v3_0/freq_div_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vssa1 0.40fF
C1231 top_pll_v3_0/s_1_n vssa1 -2.04fF
C1232 top_pll_v3_0/out_div vssa1 3.58fF
C1233 top_pll_v3_0/clk_d vssa1 1.27fF
C1234 gpio_noesd[9] vssa1 196.62fF
C1235 top_pll_v3_0/freq_div_0/inverter_min_x4_0/in vssa1 2.71fF
C1236 top_pll_v3_0/clk_5 vssa1 -0.22fF
C1237 top_pll_v3_0/clk_out_mux21 vssa1 3.89fF
C1238 top_pll_v3_0/clk_pre vssa1 1.69fF
C1239 top_pll_v3_0/freq_div_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1240 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/CLK vssa1 0.31fF
C1241 top_pll_v3_0/freq_div_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1242 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/nCLK vssa1 1.03fF
C1243 top_pll_v3_0/clk_2_f vssa1 3.30fF
C1244 top_pll_v3_0/freq_div_0/div_by_2_0/o1 vssa1 2.08fF
C1245 top_pll_v3_0/freq_div_0/div_by_2_0/nCLK_2 vssa1 1.04fF
C1246 top_pll_v3_0/freq_div_0/div_by_2_0/o2 vssa1 2.08fF
C1247 top_pll_v3_0/freq_div_0/div_by_2_0/out_div vssa1 -0.82fF
C1248 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C1249 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C1250 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C1251 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C1252 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1253 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C1254 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1255 top_pll_v3_0/freq_div_0/div_by_2_0/nout_div vssa1 2.62fF
C1256 top_pll_v3_0/freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C1257 io_analog[7] vssa1 24.25fF
C1258 top_pll_v3_0/buffer_salida_0/a_3996_n100# vssa1 48.23fF
C1259 top_pll_v3_0/buffer_salida_0/a_678_n100# vssa1 13.21fF
C1260 top_pll_v3_0/lf_vc vssa1 -60.88fF
C1261 top_pll_v3_0/loop_filter_v2_0/res_loop_filter_2/out vssa1 7.90fF
C1262 gpio_noesd[8] vssa1 303.23fF
C1263 top_pll_v3_0/loop_filter_v2_0/cap3_loop_filter_0/in vssa1 -12.03fF
C1264 top_pll_v3_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1265 top_pll_v3_0/div_by_2_0/DFlipFlop_0/CLK vssa1 0.31fF
C1266 top_pll_v3_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1267 top_pll_v3_0/div_by_2_0/DFlipFlop_0/nCLK vssa1 1.03fF
C1268 top_pll_v3_0/out_buffer_div_2 vssa1 1.57fF
C1269 top_pll_v3_0/n_out_buffer_div_2 vssa1 1.57fF
C1270 top_pll_v3_0/out_div_2 vssa1 -0.70fF
C1271 top_pll_v3_0/div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C1272 top_pll_v3_0/div_by_2_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C1273 top_pll_v3_0/div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C1274 top_pll_v3_0/div_by_2_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C1275 top_pll_v3_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1276 top_pll_v3_0/div_by_2_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C1277 top_pll_v3_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1278 top_pll_v3_0/n_out_div_2 vssa1 2.11fF
C1279 top_pll_v3_0/div_by_2_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C1280 top_pll_v3_0/nswitch vssa1 4.61fF
C1281 top_pll_v3_0/biasp vssa1 5.45fF
C1282 bias_0/iref_0 vssa1 -81.72fF
C1283 top_pll_v3_0/vco_vctrl vssa1 -30.71fF
C1284 top_pll_v3_0/pswitch vssa1 2.72fF
C1285 bias_0/iref_6 vssa1 -645.65fF
C1286 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/in vssa1 -32.98fF
C1287 io_analog[1] vssa1 73.96fF
C1288 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_1/m1_460_n1129# vssa1 1.29fF
C1289 bias_0/iref_5 vssa1 -623.45fF
C1290 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_0/in vssa1 -32.98fF
C1291 io_analog[0] vssa1 -155.24fF
C1292 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_nmos_0/m1_460_n1129# vssa1 1.29fF
C1293 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_pmos_1/m1_957_828# vssa1 -35.44fF
C1294 bias_0/iref_8 vssa1 -189.06fF
C1295 res_amp_top_0/source_follower_buff_diff_0/source_follower_buff_pmos_0/m1_957_828# vssa1 -35.44fF
C1296 bias_0/iref_7 vssa1 -205.18fF
C1297 res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_511_801# vssa1 -1.87fF
C1298 res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1384_n363# vssa1 0.47fF
C1299 gpio_noesd[5] vssa1 122.09fF
C1300 res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_448_n363# vssa1 -1.10fF
C1301 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vctrl vssa1 -2.03fF
C1302 res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_1996_n363# vssa1 -2.23fF
C1303 gpio_noesd[6] vssa1 325.91fF
C1304 gpio_noesd[4] vssa1 116.78fF
C1305 res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_964_n363# vssa1 -1.03fF
C1306 res_amp_top_0/res_amp_lin_prog_0/iref_ctrl_res_amp_0/m1_n356_n363# vssa1 0.51fF
C1307 bias_0/iref_9 vssa1 -181.57fF
C1308 res_amp_top_0/res_amp_lin_prog_0/outn vssa1 1.55fF
C1309 io_analog[3] vssa1 -119.52fF
C1310 res_amp_top_0/res_amp_lin_prog_0/outp vssa1 -4.89fF
C1311 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/vp vssa1 -4.89fF
C1312 io_analog[2] vssa1 -131.04fF
C1313 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/a_3747_261# vssa1 -0.95fF
C1314 res_amp_top_0/res_amp_lin_prog_0/outn_cap vssa1 -0.01fF
C1315 res_amp_top_0/res_amp_lin_prog_0/inverter_min_x4_0/out vssa1 4.60fF
C1316 res_amp_top_0/res_amp_lin_prog_0/res_amp_lin_0/clk vssa1 4.27fF
C1317 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_7/in vssa1 1.07fF
C1318 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinA vssa1 -0.04fF
C1319 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_7/inverter_min_1/in vssa1 1.03fF
C1320 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_6/inverter_min_1/in vssa1 1.03fF
C1321 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_5/in vssa1 1.07fF
C1322 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_5/inverter_min_1/in vssa1 1.03fF
C1323 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_4/inverter_min_1/in vssa1 1.03fF
C1324 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_3/in vssa1 1.07fF
C1325 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_3/inverter_min_1/in vssa1 1.03fF
C1326 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_1/in vssa1 1.07fF
C1327 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_1/inverter_min_1/in vssa1 1.03fF
C1328 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_2/inverter_min_1/in vssa1 1.03fF
C1329 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_0/inverter_min_1/in vssa1 1.03fF
C1330 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/in vssa1 1.07fF
C1331 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinB vssa1 -7.88fF
C1332 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_13/inverter_min_1/in vssa1 1.03fF
C1333 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_12/inverter_min_1/in vssa1 1.03fF
C1334 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_11/in vssa1 1.07fF
C1335 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_11/inverter_min_1/in vssa1 1.03fF
C1336 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/m1_21_n341# vssa1 0.72fF
C1337 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_10/inverter_min_1/in vssa1 1.03fF
C1338 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/nand_logic_0/in1 vssa1 1.54fF
C1339 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_6/sel_b vssa1 2.03fF
C1340 gpio_noesd[3] vssa1 213.06fF
C1341 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_5/out vssa1 -1.67fF
C1342 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_5/sel_b vssa1 2.03fF
C1343 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/DinA vssa1 -2.58fF
C1344 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/out vssa1 -2.25fF
C1345 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_4/sel_b vssa1 2.03fF
C1346 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/out vssa1 -2.69fF
C1347 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/DinB vssa1 -4.96fF
C1348 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_3/sel_b vssa1 2.03fF
C1349 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/out vssa1 -4.71fF
C1350 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_2/sel_b vssa1 2.03fF
C1351 gpio_noesd[2] vssa1 216.13fF
C1352 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/DinA vssa1 0.63fF
C1353 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/out vssa1 -2.49fF
C1354 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/DinB vssa1 -3.92fF
C1355 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_1/sel_b vssa1 2.03fF
C1356 gpio_noesd[1] vssa1 230.09fF
C1357 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/out vssa1 -0.27fF
C1358 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/DinB vssa1 -0.97fF
C1359 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/mux_2to1_logic_0/sel_b vssa1 2.03fF
C1360 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_9/in vssa1 1.07fF
C1361 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_9/inverter_min_1/in vssa1 1.03fF
C1362 res_amp_top_0/res_amp_lin_prog_0/delay_cell_buff_0/buffer_no_inv_x05_8/inverter_min_1/in vssa1 1.03fF
C1363 res_amp_top_0/res_amp_lin_prog_0/outp_cap vssa1 -7.66fF
C1364 res_amp_top_0/res_amp_sync_v2_0/nand_logic_1/m1_21_n341# vssa1 0.72fF
C1365 res_amp_top_0/res_amp_sync_v2_0/nand_logic_0/m1_21_n341# vssa1 0.72fF
C1366 res_amp_top_0/res_amp_lin_prog_0/clk vssa1 -8.26fF
C1367 res_amp_top_0/res_amp_sync_v2_0/inverter_min_x4_4/out vssa1 5.85fF
C1368 res_amp_top_0/res_amp_sync_v2_0/rst vssa1 -7.88fF
C1369 res_amp_top_0/res_amp_sync_v2_0/nand_logic_1/out vssa1 1.70fF
C1370 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/Q vssa1 -2.08fF
C1371 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/m1_657_280# vssa1 0.57fF
C1372 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/nQ vssa1 0.48fF
C1373 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/D vssa1 -1.73fF
C1374 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/latch_diff_0/m1_657_280# vssa1 0.57fF
C1375 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/latch_diff_1/nD vssa1 0.57fF
C1376 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1377 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/latch_diff_0/D vssa1 0.96fF
C1378 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1379 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/D vssa1 1.83fF
C1380 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_4/latch_diff_0/nD vssa1 1.14fF
C1381 res_amp_top_0/res_amp_sync_v2_0/nand_logic_0/out vssa1 1.20fF
C1382 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/Q vssa1 -2.94fF
C1383 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/m1_657_280# vssa1 0.57fF
C1384 io_analog[4] vssa1 -253.69fF
C1385 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/nQ vssa1 0.48fF
C1386 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/D vssa1 -1.73fF
C1387 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/latch_diff_0/m1_657_280# vssa1 0.57fF
C1388 io_analog[6] vssa1 -26.69fF
C1389 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/latch_diff_1/nD vssa1 0.57fF
C1390 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1391 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/latch_diff_0/D vssa1 0.96fF
C1392 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1393 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/D vssa1 0.79fF
C1394 vdda1 vssa1 7499.69fF
C1395 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_3/latch_diff_0/nD vssa1 1.14fF
C1396 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/Q vssa1 -1.08fF
C1397 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/latch_diff_1/m1_657_280# vssa1 0.57fF
C1398 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/nQ vssa1 0.48fF
C1399 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/latch_diff_1/D vssa1 -1.73fF
C1400 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/latch_diff_0/m1_657_280# vssa1 0.57fF
C1401 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/latch_diff_1/nD vssa1 0.57fF
C1402 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1403 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/latch_diff_0/D vssa1 0.96fF
C1404 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1405 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/D vssa1 -0.38fF
C1406 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_2/latch_diff_0/nD vssa1 1.14fF
C1407 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/latch_diff_1/m1_657_280# vssa1 0.57fF
C1408 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/nQ vssa1 0.48fF
C1409 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/latch_diff_1/D vssa1 -1.73fF
C1410 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/latch_diff_0/m1_657_280# vssa1 0.57fF
C1411 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/latch_diff_1/nD vssa1 0.57fF
C1412 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1413 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/latch_diff_0/D vssa1 0.96fF
C1414 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1415 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/D vssa1 -1.04fF
C1416 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_1/latch_diff_0/nD vssa1 1.14fF
C1417 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/Q vssa1 -4.73fF
C1418 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C1419 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/nQ vssa1 0.48fF
C1420 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C1421 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C1422 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C1423 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1424 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C1425 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1426 res_amp_top_0/res_amp_sync_v2_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
.ends

