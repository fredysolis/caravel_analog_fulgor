**.subckt tb_div_by_5_pex_c
VSS vss GND {vss} 
VDD vdd vss {vdd} 
x1 nclk_2 vss A vdd clk_2 net14 net15 net16 net17 div_by_2_pex_c
Vref net1 vss PULSE(0 {vin} 0 1p 1p {Tref/2} {Tref}) DC {vin} AC 0 
x3 vdd net2 net1 vss inverter_min_x2_pex_c
x4 vdd A net2 vss inverter_min_x4_pex_c
x5 vss vdd net10 net11 clk_5 net9 net8 PFD_pex_c
x2 vdd clk_5 clk_2_buf vss nclk_2_buf net3 net4 net6 net7 net5 div_by_5_pex_c
x6 vdd net12 clk_2 vss inverter_min_x2_pex_c
x7 vdd clk_2_buf net12 vss inverter_min_x4_pex_c
x8 vdd net13 nclk_2 vss inverter_min_x2_pex_c
x9 vdd nclk_2_buf net13 vss inverter_min_x4_pex_c
**** begin user architecture code



* Parameters
.param kp = 1.0
.param vdd = kp*1.8
.param vss = 0.0
.param vin = vdd
.param fref = 1e9
.param Tref = 1/fref
.param C = 1f
.param iref=100u

.options TEMP = 100.0
.options RSHUNT = 1e20

* Models
.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib SS
.include ~/caravel_analog_fulgor/xschem/simulations/inverter_min_x2_pex_c.spice
.include ~/caravel_analog_fulgor/xschem/simulations/inverter_min_x4_pex_c.spice
.include ~/caravel_analog_fulgor/xschem/simulations/div_by_2_pex_c.spice
.include ~/caravel_analog_fulgor/xschem/simulations/div_by_5_pex_c.spice
.include ~/caravel_analog_fulgor/xschem/simulations/PFD_pex_c.spice

* Data to save
.save all

.ic v(A) = 0.0
.ic v(x2.q0) = 0.0
.ic v(x2.nq0) = 0.0
.ic v(x2.q1) = 0.0
.ic v(x2.nq1) = 0.0
.ic v(x2.q1_shift) = 0.0
.ic v(x2.nq1_shift) = 0.0
.ic v(x2.q2) = 0.0
.ic v(x2.nq2) = 0.0
.ic v(x2.x1.a) = 0.0
.ic v(x2.x1.na) = 0.0
.ic v(x2.x1.D_d) = 0.0
.ic v(x2.x1.nD_d) = 0.0
.ic v(clk_2) = 0.0
.ic v(nclk_2) = 0.0
.ic v(clk_5)

* Simulation
.control
	tran 0.01ns 200ns
	write tb_div_by_5_tran.raw
	plot v(clk_2) v(A) v(nclk_2)+2 v(A)+2
	plot v(clk_5) v(clk_2_buf) v(A)
.endc



**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
