magic
tech sky130A
magscale 1 2
timestamp 1623948030
<< nwell >>
rect 2984 2989 4228 3068
rect 3203 118 4219 142
rect 3203 84 4228 118
rect 3203 83 4219 84
rect 3203 79 4228 83
rect 2984 0 4228 79
<< pwell >>
rect 2983 1339 4228 1819
<< locali >>
rect 1986 2123 2002 2157
rect 2224 2123 2240 2157
<< metal1 >>
rect 2984 3022 4228 3038
rect 2947 2998 4228 3022
rect -1244 2957 4228 2998
rect -1244 2944 3720 2957
rect 2947 2931 3720 2944
rect 2986 2918 3533 2931
rect -190 2228 -180 2356
rect -116 2228 -106 2356
rect 2984 2267 2994 2323
rect 3218 2267 3228 2323
rect 3352 2253 3753 2333
rect 4061 2249 4228 2327
rect 1990 2121 2000 2173
rect 2226 2121 2236 2173
rect 1990 2117 2236 2121
rect 2915 1848 2984 1864
rect 2915 1825 3020 1848
rect 2915 1730 4224 1825
rect 2915 1700 4228 1730
rect -1244 1498 1313 1570
rect 2915 1369 3020 1700
rect 3412 1369 3726 1700
rect 2915 1339 4228 1369
rect 2915 1321 3726 1339
rect 2915 1282 3556 1321
rect 2915 1266 3130 1282
rect 2915 1246 3020 1266
rect 2915 1204 2984 1246
rect 1992 947 2238 951
rect 1992 895 2002 947
rect 2228 895 2238 947
rect -150 712 -140 840
rect -76 712 -66 840
rect 2981 748 2991 804
rect 3215 748 3225 804
rect 3352 736 3753 816
rect 4061 742 4228 820
rect 2915 148 4220 164
rect 2915 30 4228 148
<< via1 >>
rect -180 2228 -116 2356
rect 2994 2267 3218 2323
rect 2000 2121 2226 2173
rect 2002 895 2228 947
rect -140 712 -76 840
rect 2991 748 3215 804
<< metal2 >>
rect -180 2356 -116 2366
rect -180 2218 -116 2228
rect 2081 2321 2145 2331
rect 2000 2173 2081 2183
rect 2994 2323 3218 2333
rect 2994 2257 3218 2267
rect 2145 2173 2226 2183
rect 2000 2111 2226 2121
rect 250 1569 306 1579
rect 2555 1570 2611 1580
rect 306 1477 2555 1549
rect 306 1475 323 1477
rect 250 1447 306 1457
rect 2611 1477 2621 1549
rect 2555 1448 2611 1458
rect 2002 947 2228 957
rect 2002 885 2083 895
rect -140 840 -76 850
rect 2147 885 2228 895
rect 2083 734 2147 744
rect 2991 804 3215 814
rect 2991 738 3215 748
rect -140 702 -76 712
<< via2 >>
rect -180 2228 -116 2356
rect 2081 2173 2145 2321
rect 2994 2267 3218 2323
rect 2081 2121 2145 2173
rect 250 1457 306 1569
rect 2555 1458 2611 1570
rect 2083 895 2147 900
rect -140 712 -76 840
rect 2083 744 2147 895
rect 2991 748 3215 804
<< metal3 >>
rect -190 2356 -106 2361
rect -997 804 -937 2264
rect -190 2228 -180 2356
rect -116 2228 -106 2356
rect -190 2223 -106 2228
rect 2071 2321 2155 2326
rect 2071 2121 2081 2321
rect 2145 2121 2155 2321
rect 2763 2325 2823 2474
rect 2984 2325 3228 2328
rect 2763 2323 3246 2325
rect 2763 2267 2994 2323
rect 3218 2267 3246 2323
rect 2763 2265 3246 2267
rect 2071 2116 2155 2121
rect 2553 1575 2613 2258
rect 240 1569 316 1574
rect 240 1457 250 1569
rect 306 1457 316 1569
rect 240 1452 316 1457
rect 2545 1570 2621 1575
rect 2545 1458 2555 1570
rect 2611 1458 2621 1570
rect 2545 1453 2621 1458
rect 2073 945 2157 950
rect -150 840 -66 845
rect -150 712 -140 840
rect -76 712 -66 840
rect 2073 744 2083 945
rect 2147 744 2157 945
rect 2073 739 2157 744
rect -150 707 -66 712
rect 2553 596 2613 1453
rect 2763 810 2823 2265
rect 2984 2262 3228 2265
rect 2981 808 3225 809
rect 2977 804 3225 808
rect 2977 748 2991 804
rect 3215 748 3225 804
rect 2977 743 3225 748
rect 2977 596 3037 743
rect 2528 536 3037 596
<< via3 >>
rect -180 2228 -116 2356
rect 2081 2121 2145 2321
rect -140 712 -76 840
rect 2083 900 2147 945
rect 2083 744 2147 900
<< metal4 >>
rect -181 2356 -115 2357
rect -181 2228 -180 2356
rect -116 2324 -115 2356
rect -116 2322 2139 2324
rect -116 2321 2146 2322
rect -116 2260 2081 2321
rect -116 2228 -115 2260
rect -181 2227 -115 2228
rect 2080 2121 2081 2260
rect 2145 2121 2146 2321
rect 2080 2120 2146 2121
rect 2082 945 2148 946
rect -141 840 -75 841
rect -141 712 -140 840
rect -76 808 -75 840
rect 2082 808 2083 945
rect -76 744 2083 808
rect 2147 744 2148 945
rect -76 712 -75 744
rect 2082 743 2148 744
rect -141 711 -75 712
use DFlipFlop  DFlipFlop_0
timestamp 1623898709
transform 1 0 1244 0 -1 3068
box -1244 0 1740 3068
use clock_inverter  clock_inverter_0
timestamp 1623799048
transform 1 0 -1244 0 1 0
box 0 0 1244 3068
use inverter_min_x2  inverter_min_x2_0
timestamp 1623898709
transform 1 0 3037 0 -1 723
box -53 -615 473 655
use inverter_min_x2  inverter_min_x2_1
timestamp 1623898709
transform 1 0 3037 0 1 2345
box -53 -615 473 655
use inverter_min_x4  inverter_min_x4_0
timestamp 1623895985
transform 1 0 3563 0 1 2346
box -53 -616 665 643
use inverter_min_x4  inverter_min_x4_1
timestamp 1623895985
transform 1 0 3563 0 -1 723
box -53 -616 665 643
<< labels >>
rlabel metal1 -1244 2944 2984 2998 1 vdd
rlabel metal1 -1244 1498 1313 1570 1 vss
rlabel metal3 -997 1498 -937 1570 1 CLK
rlabel metal3 2553 1570 2613 2258 1 nout_div
rlabel metal3 2763 810 2823 2474 1 out_div
rlabel metal1 4061 2249 4228 2327 1 CLK_2
rlabel metal1 3352 2253 3753 2333 1 o1
rlabel metal1 3352 736 3753 816 1 o2
rlabel metal1 4061 742 4228 820 1 nCLK_2
<< end >>
