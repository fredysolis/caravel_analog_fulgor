magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< pwell >>
rect -1367 -285 1367 285
<< nmos >>
rect -1167 -75 -1137 75
rect -1071 -75 -1041 75
rect -975 -75 -945 75
rect -879 -75 -849 75
rect -783 -75 -753 75
rect -687 -75 -657 75
rect -591 -75 -561 75
rect -495 -75 -465 75
rect -399 -75 -369 75
rect -303 -75 -273 75
rect -207 -75 -177 75
rect -111 -75 -81 75
rect -15 -75 15 75
rect 81 -75 111 75
rect 177 -75 207 75
rect 273 -75 303 75
rect 369 -75 399 75
rect 465 -75 495 75
rect 561 -75 591 75
rect 657 -75 687 75
rect 753 -75 783 75
rect 849 -75 879 75
rect 945 -75 975 75
rect 1041 -75 1071 75
rect 1137 -75 1167 75
<< ndiff >>
rect -1229 63 -1167 75
rect -1229 -63 -1217 63
rect -1183 -63 -1167 63
rect -1229 -75 -1167 -63
rect -1137 63 -1071 75
rect -1137 -63 -1121 63
rect -1087 -63 -1071 63
rect -1137 -75 -1071 -63
rect -1041 63 -975 75
rect -1041 -63 -1025 63
rect -991 -63 -975 63
rect -1041 -75 -975 -63
rect -945 63 -879 75
rect -945 -63 -929 63
rect -895 -63 -879 63
rect -945 -75 -879 -63
rect -849 63 -783 75
rect -849 -63 -833 63
rect -799 -63 -783 63
rect -849 -75 -783 -63
rect -753 63 -687 75
rect -753 -63 -737 63
rect -703 -63 -687 63
rect -753 -75 -687 -63
rect -657 63 -591 75
rect -657 -63 -641 63
rect -607 -63 -591 63
rect -657 -75 -591 -63
rect -561 63 -495 75
rect -561 -63 -545 63
rect -511 -63 -495 63
rect -561 -75 -495 -63
rect -465 63 -399 75
rect -465 -63 -449 63
rect -415 -63 -399 63
rect -465 -75 -399 -63
rect -369 63 -303 75
rect -369 -63 -353 63
rect -319 -63 -303 63
rect -369 -75 -303 -63
rect -273 63 -207 75
rect -273 -63 -257 63
rect -223 -63 -207 63
rect -273 -75 -207 -63
rect -177 63 -111 75
rect -177 -63 -161 63
rect -127 -63 -111 63
rect -177 -75 -111 -63
rect -81 63 -15 75
rect -81 -63 -65 63
rect -31 -63 -15 63
rect -81 -75 -15 -63
rect 15 63 81 75
rect 15 -63 31 63
rect 65 -63 81 63
rect 15 -75 81 -63
rect 111 63 177 75
rect 111 -63 127 63
rect 161 -63 177 63
rect 111 -75 177 -63
rect 207 63 273 75
rect 207 -63 223 63
rect 257 -63 273 63
rect 207 -75 273 -63
rect 303 63 369 75
rect 303 -63 319 63
rect 353 -63 369 63
rect 303 -75 369 -63
rect 399 63 465 75
rect 399 -63 415 63
rect 449 -63 465 63
rect 399 -75 465 -63
rect 495 63 561 75
rect 495 -63 511 63
rect 545 -63 561 63
rect 495 -75 561 -63
rect 591 63 657 75
rect 591 -63 607 63
rect 641 -63 657 63
rect 591 -75 657 -63
rect 687 63 753 75
rect 687 -63 703 63
rect 737 -63 753 63
rect 687 -75 753 -63
rect 783 63 849 75
rect 783 -63 799 63
rect 833 -63 849 63
rect 783 -75 849 -63
rect 879 63 945 75
rect 879 -63 895 63
rect 929 -63 945 63
rect 879 -75 945 -63
rect 975 63 1041 75
rect 975 -63 991 63
rect 1025 -63 1041 63
rect 975 -75 1041 -63
rect 1071 63 1137 75
rect 1071 -63 1087 63
rect 1121 -63 1137 63
rect 1071 -75 1137 -63
rect 1167 63 1229 75
rect 1167 -63 1183 63
rect 1217 -63 1229 63
rect 1167 -75 1229 -63
<< ndiffc >>
rect -1217 -63 -1183 63
rect -1121 -63 -1087 63
rect -1025 -63 -991 63
rect -929 -63 -895 63
rect -833 -63 -799 63
rect -737 -63 -703 63
rect -641 -63 -607 63
rect -545 -63 -511 63
rect -449 -63 -415 63
rect -353 -63 -319 63
rect -257 -63 -223 63
rect -161 -63 -127 63
rect -65 -63 -31 63
rect 31 -63 65 63
rect 127 -63 161 63
rect 223 -63 257 63
rect 319 -63 353 63
rect 415 -63 449 63
rect 511 -63 545 63
rect 607 -63 641 63
rect 703 -63 737 63
rect 799 -63 833 63
rect 895 -63 929 63
rect 991 -63 1025 63
rect 1087 -63 1121 63
rect 1183 -63 1217 63
<< psubdiff >>
rect 1297 153 1331 215
rect 1297 -215 1331 -153
rect -1297 -249 -1235 -215
rect 1235 -249 1331 -215
<< psubdiffcont >>
rect 1297 -153 1331 153
rect -1235 -249 1235 -215
<< poly >>
rect -1167 101 1167 167
rect -1167 75 -1137 101
rect -1071 75 -1041 101
rect -975 75 -945 101
rect -879 75 -849 101
rect -783 75 -753 101
rect -687 75 -657 101
rect -591 75 -561 101
rect -495 75 -465 101
rect -399 75 -369 101
rect -303 75 -273 101
rect -207 75 -177 101
rect -111 75 -81 101
rect -15 75 15 101
rect 81 75 111 101
rect 177 75 207 101
rect 273 75 303 101
rect 369 75 399 101
rect 465 75 495 101
rect 561 75 591 101
rect 657 75 687 101
rect 753 75 783 101
rect 849 75 879 101
rect 945 75 975 101
rect 1041 75 1071 101
rect 1137 75 1167 101
rect -1167 -101 -1137 -75
rect -1071 -101 -1041 -75
rect -975 -101 -945 -75
rect -879 -101 -849 -75
rect -783 -101 -753 -75
rect -687 -101 -657 -75
rect -591 -101 -561 -75
rect -495 -101 -465 -75
rect -399 -101 -369 -75
rect -303 -101 -273 -75
rect -207 -101 -177 -75
rect -111 -101 -81 -75
rect -15 -101 15 -75
rect 81 -101 111 -75
rect 177 -101 207 -75
rect 273 -101 303 -75
rect 369 -101 399 -75
rect 465 -101 495 -75
rect 561 -101 591 -75
rect 657 -101 687 -75
rect 753 -101 783 -75
rect 849 -101 879 -75
rect 945 -101 975 -75
rect 1041 -101 1071 -75
rect 1137 -101 1167 -75
<< locali >>
rect 1297 153 1331 215
rect -1217 63 -1183 79
rect -1217 -79 -1183 -63
rect -1121 63 -1087 79
rect -1121 -79 -1087 -63
rect -1025 63 -991 79
rect -1025 -79 -991 -63
rect -929 63 -895 79
rect -929 -79 -895 -63
rect -833 63 -799 79
rect -833 -79 -799 -63
rect -737 63 -703 79
rect -737 -79 -703 -63
rect -641 63 -607 79
rect -641 -79 -607 -63
rect -545 63 -511 79
rect -545 -79 -511 -63
rect -449 63 -415 79
rect -449 -79 -415 -63
rect -353 63 -319 79
rect -353 -79 -319 -63
rect -257 63 -223 79
rect -257 -79 -223 -63
rect -161 63 -127 79
rect -161 -79 -127 -63
rect -65 63 -31 79
rect -65 -79 -31 -63
rect 31 63 65 79
rect 31 -79 65 -63
rect 127 63 161 79
rect 127 -79 161 -63
rect 223 63 257 79
rect 223 -79 257 -63
rect 319 63 353 79
rect 319 -79 353 -63
rect 415 63 449 79
rect 415 -79 449 -63
rect 511 63 545 79
rect 511 -79 545 -63
rect 607 63 641 79
rect 607 -79 641 -63
rect 703 63 737 79
rect 703 -79 737 -63
rect 799 63 833 79
rect 799 -79 833 -63
rect 895 63 929 79
rect 895 -79 929 -63
rect 991 63 1025 79
rect 991 -79 1025 -63
rect 1087 63 1121 79
rect 1087 -79 1121 -63
rect 1183 63 1217 79
rect 1183 -79 1217 -63
rect 1297 -215 1331 -153
rect -1297 -249 -1235 -215
rect 1235 -249 1331 -215
<< viali >>
rect -1217 -63 -1183 63
rect -1121 -63 -1087 63
rect -1025 -63 -991 63
rect -929 -63 -895 63
rect -833 -63 -799 63
rect -737 -63 -703 63
rect -641 -63 -607 63
rect -545 -63 -511 63
rect -449 -63 -415 63
rect -353 -63 -319 63
rect -257 -63 -223 63
rect -161 -63 -127 63
rect -65 -63 -31 63
rect 31 -63 65 63
rect 127 -63 161 63
rect 223 -63 257 63
rect 319 -63 353 63
rect 415 -63 449 63
rect 511 -63 545 63
rect 607 -63 641 63
rect 703 -63 737 63
rect 799 -63 833 63
rect 895 -63 929 63
rect 991 -63 1025 63
rect 1087 -63 1121 63
rect 1183 -63 1217 63
<< metal1 >>
rect -1223 63 -1177 75
rect -1223 -63 -1217 63
rect -1183 -63 -1177 63
rect -1223 -75 -1177 -63
rect -1127 63 -1081 75
rect -1127 -63 -1121 63
rect -1087 -63 -1081 63
rect -1127 -75 -1081 -63
rect -1031 63 -985 75
rect -1031 -63 -1025 63
rect -991 -63 -985 63
rect -1031 -75 -985 -63
rect -935 63 -889 75
rect -935 -63 -929 63
rect -895 -63 -889 63
rect -935 -75 -889 -63
rect -839 63 -793 75
rect -839 -63 -833 63
rect -799 -63 -793 63
rect -839 -75 -793 -63
rect -743 63 -697 75
rect -743 -63 -737 63
rect -703 -63 -697 63
rect -743 -75 -697 -63
rect -647 63 -601 75
rect -647 -63 -641 63
rect -607 -63 -601 63
rect -647 -75 -601 -63
rect -551 63 -505 75
rect -551 -63 -545 63
rect -511 -63 -505 63
rect -551 -75 -505 -63
rect -455 63 -409 75
rect -455 -63 -449 63
rect -415 -63 -409 63
rect -455 -75 -409 -63
rect -359 63 -313 75
rect -359 -63 -353 63
rect -319 -63 -313 63
rect -359 -75 -313 -63
rect -263 63 -217 75
rect -263 -63 -257 63
rect -223 -63 -217 63
rect -263 -75 -217 -63
rect -167 63 -121 75
rect -167 -63 -161 63
rect -127 -63 -121 63
rect -167 -75 -121 -63
rect -71 63 -25 75
rect -71 -63 -65 63
rect -31 -63 -25 63
rect -71 -75 -25 -63
rect 25 63 71 75
rect 25 -63 31 63
rect 65 -63 71 63
rect 25 -75 71 -63
rect 121 63 167 75
rect 121 -63 127 63
rect 161 -63 167 63
rect 121 -75 167 -63
rect 217 63 263 75
rect 217 -63 223 63
rect 257 -63 263 63
rect 217 -75 263 -63
rect 313 63 359 75
rect 313 -63 319 63
rect 353 -63 359 63
rect 313 -75 359 -63
rect 409 63 455 75
rect 409 -63 415 63
rect 449 -63 455 63
rect 409 -75 455 -63
rect 505 63 551 75
rect 505 -63 511 63
rect 545 -63 551 63
rect 505 -75 551 -63
rect 601 63 647 75
rect 601 -63 607 63
rect 641 -63 647 63
rect 601 -75 647 -63
rect 697 63 743 75
rect 697 -63 703 63
rect 737 -63 743 63
rect 697 -75 743 -63
rect 793 63 839 75
rect 793 -63 799 63
rect 833 -63 839 63
rect 793 -75 839 -63
rect 889 63 935 75
rect 889 -63 895 63
rect 929 -63 935 63
rect 889 -75 935 -63
rect 985 63 1031 75
rect 985 -63 991 63
rect 1025 -63 1031 63
rect 985 -75 1031 -63
rect 1081 63 1127 75
rect 1081 -63 1087 63
rect 1121 -63 1127 63
rect 1081 -75 1127 -63
rect 1177 63 1223 75
rect 1177 -63 1183 63
rect 1217 -63 1223 63
rect 1177 -75 1223 -63
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1314 -232 1314 232
string parameters w 0.75 l 0.150 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
