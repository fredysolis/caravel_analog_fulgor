magic
tech sky130A
magscale 1 2
timestamp 1623450397
<< nwell >>
rect -263 -309 263 309
<< pmos >>
rect -63 -90 -33 90
rect 33 -90 63 90
<< pdiff >>
rect -125 78 -63 90
rect -125 -78 -113 78
rect -79 -78 -63 78
rect -125 -90 -63 -78
rect -33 78 33 90
rect -33 -78 -17 78
rect 17 -78 33 78
rect -33 -90 33 -78
rect 63 78 125 90
rect 63 -78 79 78
rect 113 -78 125 78
rect 63 -90 125 -78
<< pdiffc >>
rect -113 -78 -79 78
rect -17 -78 17 78
rect 79 -78 113 78
<< nsubdiff >>
rect -193 239 -131 273
rect 131 239 193 273
<< nsubdiffcont >>
rect -131 239 131 273
<< poly >>
rect -63 90 -33 116
rect 33 90 63 116
rect -63 -121 -33 -90
rect -99 -187 -33 -121
rect 33 -121 63 -90
rect 33 -187 99 -121
<< locali >>
rect -193 239 -131 273
rect 131 239 193 273
rect -113 78 -79 94
rect -113 -94 -79 -78
rect -17 78 17 94
rect -17 -94 17 -78
rect 79 78 113 94
rect 79 -94 113 -78
<< viali >>
rect -113 -78 -79 78
rect -17 -78 17 78
rect 79 -78 113 78
<< metal1 >>
rect -119 78 -73 90
rect -119 -78 -113 78
rect -79 -78 -73 78
rect -119 -90 -73 -78
rect -23 78 23 90
rect -23 -78 -17 78
rect 17 -78 23 78
rect -23 -90 23 -78
rect 73 78 119 90
rect 73 -78 79 78
rect 113 -78 119 78
rect 73 -90 119 -78
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -210 -256 210 256
string parameters w 0.9 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
