magic
tech sky130A
magscale 1 2
timestamp 1624064496
<< nwell >>
rect -363 387 931 1955
<< pwell >>
rect -363 -680 931 387
rect -363 -771 162 -680
rect 184 -771 931 -680
rect -363 -1002 931 -771
<< psubdiff >>
rect 608 -174 632 -140
rect 790 -174 814 -140
rect -255 -966 -231 -932
rect 799 -966 823 -932
<< nsubdiff >>
rect -247 1871 -223 1905
rect 807 1871 831 1905
<< psubdiffcont >>
rect 632 -174 790 -140
rect -231 -966 799 -932
<< nsubdiffcont >>
rect -223 1871 807 1905
<< locali >>
rect -239 1871 -223 1905
rect 807 1871 823 1905
<< viali >>
rect -223 1871 807 1905
rect 104 1742 454 1776
rect 104 1214 138 1742
rect 420 1214 454 1742
rect 104 1180 454 1214
rect 536 -85 886 -51
rect 536 -174 632 -140
rect 632 -174 790 -140
rect 790 -174 886 -140
rect 106 -285 456 -251
rect 106 -796 140 -285
rect 422 -796 456 -285
rect 106 -837 459 -796
rect -327 -966 -231 -932
rect -231 -966 799 -932
rect 799 -966 895 -932
<< metal1 >>
rect -363 1905 931 1911
rect -363 1871 -223 1905
rect 807 1871 931 1905
rect -363 1776 931 1871
rect -363 1736 104 1776
rect 68 1180 104 1736
rect 138 1736 420 1742
rect 138 1220 144 1736
rect 185 1641 195 1699
rect 307 1641 317 1699
rect 247 1630 311 1641
rect 347 1595 420 1736
rect 174 1278 184 1569
rect 252 1278 262 1569
rect 342 1291 420 1595
rect 414 1220 420 1291
rect 138 1214 420 1220
rect 454 1736 931 1776
rect 454 1180 500 1736
rect 68 1108 500 1180
rect 209 897 261 907
rect 209 607 261 617
rect 68 361 78 413
rect 286 361 296 413
rect 356 361 366 413
rect 490 361 500 413
rect 631 361 641 413
rect 693 361 703 413
rect 209 167 261 177
rect 644 173 690 361
rect 760 89 770 234
rect 831 89 841 234
rect 209 27 261 37
rect 619 8 629 60
rect 733 8 743 60
rect 61 -174 81 -45
rect 500 -51 931 -45
rect 500 -85 536 -51
rect 886 -85 931 -51
rect 500 -140 931 -85
rect 500 -174 536 -140
rect 886 -174 931 -140
rect 61 -220 931 -174
rect 61 -251 932 -220
rect 61 -790 106 -251
rect 456 -256 932 -251
rect 456 -257 737 -256
rect -363 -837 106 -790
rect 140 -291 422 -285
rect 140 -790 146 -291
rect 416 -364 422 -291
rect 191 -651 201 -374
rect 258 -651 268 -374
rect 249 -701 313 -692
rect 178 -704 313 -701
rect 178 -756 184 -704
rect 308 -756 318 -704
rect 347 -790 422 -364
rect 140 -796 422 -790
rect 456 -291 468 -257
rect 456 -790 462 -291
rect 456 -796 931 -790
rect 459 -837 931 -796
rect -363 -932 931 -837
rect -363 -966 -327 -932
rect 895 -966 931 -932
rect -363 -972 931 -966
<< via1 >>
rect 195 1641 307 1699
rect 184 1278 252 1569
rect 209 617 261 897
rect 78 361 286 413
rect 366 361 490 413
rect 641 361 693 413
rect 209 37 261 167
rect 770 89 831 234
rect 629 8 733 60
rect 201 -651 258 -374
rect 184 -756 308 -704
<< metal2 >>
rect 195 1699 307 1709
rect 80 1641 195 1682
rect 307 1641 312 1682
rect 80 1629 312 1641
rect 184 1574 252 1579
rect 184 1569 261 1574
rect 252 1278 261 1569
rect 184 1268 261 1278
rect 209 897 261 1268
rect 209 607 261 617
rect 78 413 286 423
rect 68 361 78 413
rect 78 351 286 361
rect 366 413 490 423
rect 641 413 693 423
rect 490 361 641 413
rect 693 361 931 413
rect 366 351 490 361
rect 641 351 693 361
rect 813 244 874 245
rect 770 235 874 244
rect 770 234 813 235
rect 209 167 261 177
rect 831 89 874 90
rect 770 80 874 89
rect 770 79 831 80
rect 209 -364 261 37
rect 629 62 733 72
rect 629 -4 733 6
rect 201 -374 261 -364
rect 258 -463 261 -374
rect 201 -661 258 -651
rect 184 -703 308 -694
rect 699 -703 886 -702
rect 73 -704 321 -703
rect 73 -756 184 -704
rect 308 -756 321 -704
rect 699 -713 900 -703
rect 699 -748 797 -713
rect 73 -758 321 -756
rect 184 -766 308 -758
rect 797 -781 900 -771
<< via2 >>
rect 813 234 874 235
rect 813 90 831 234
rect 831 90 874 234
rect 629 60 733 62
rect 629 8 733 60
rect 629 6 733 8
rect 797 -771 900 -713
<< metal3 >>
rect 803 239 884 240
rect 803 235 886 239
rect 803 90 813 235
rect 874 90 886 235
rect 803 85 886 90
rect 619 62 743 67
rect 619 6 629 62
rect 733 6 743 62
rect 619 1 743 6
rect 650 -194 710 1
rect 819 -708 886 85
rect 787 -713 910 -708
rect 787 -771 797 -713
rect 900 -771 910 -713
rect 787 -776 910 -771
use cap_vco  cap_vco_0
timestamp 1624049879
transform 1 0 -37 0 1 -744
box 554 -6 926 514
use sky130_fd_pr__nfet_01v8_EDT3AT  sky130_fd_pr__nfet_01v8_EDT3AT_0
timestamp 1624049879
transform 1 0 711 0 1 100
box -211 -221 211 221
use sky130_fd_pr__nfet_01v8_CBSTVW  sky130_fd_pr__nfet_01v8_CBSTVW_0
timestamp 1624058804
transform 1 0 281 0 1 -544
box -211 -329 211 329
use inverter_csvco  inverter_csvco_0
timestamp 1624049879
transform 1 0 68 0 1 387
box 0 -597 432 757
use sky130_fd_pr__pfet_01v8_MJP3BN  sky130_fd_pr__pfet_01v8_MJP3BN_0
timestamp 1624058804
transform 1 0 279 0 1 1478
box -211 -334 211 334
<< labels >>
rlabel metal2 68 361 78 413 1 in
rlabel metal3 650 -194 710 6 1 D0
rlabel metal2 693 361 931 413 1 out
rlabel metal2 73 -758 177 -703 1 vctrl
rlabel metal1 -363 1776 931 1871 1 vdd
rlabel metal1 -363 -932 931 -837 1 vss
<< end >>
