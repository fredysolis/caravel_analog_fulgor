magic
tech sky130A
magscale 1 2
timestamp 1624019461
<< metal3 >>
rect -6469 2200 -2301 6400
rect -2150 2200 2018 6400
rect 2169 6372 6468 6400
rect 2169 2228 6384 6372
rect 6448 2228 6468 6372
rect 2169 2200 6468 2228
rect -6469 -2100 -2301 2100
rect -2150 -2100 2018 2100
rect 2169 2072 6468 2100
rect 2169 -2072 6384 2072
rect 6448 -2072 6468 2072
rect 2169 -2100 6468 -2072
rect -6469 -6400 -2301 -2200
rect -2150 -6400 2018 -2200
rect 2169 -2228 6468 -2200
rect 2169 -6372 6384 -2228
rect 6448 -6372 6468 -2228
rect 2169 -6400 6468 -6372
<< via3 >>
rect 6384 2228 6448 6372
rect 6384 -2072 6448 2072
rect 6384 -6372 6448 -2228
<< mimcap >>
rect -6369 6260 -2369 6300
rect -6369 2340 -6329 6260
rect -2409 2340 -2369 6260
rect -6369 2300 -2369 2340
rect -2050 6260 1950 6300
rect -2050 2340 -2010 6260
rect 1910 2340 1950 6260
rect -2050 2300 1950 2340
rect 2269 6260 6269 6300
rect 2269 2340 2309 6260
rect 6229 2340 6269 6260
rect 2269 2300 6269 2340
rect -6369 1960 -2369 2000
rect -6369 -1960 -6329 1960
rect -2409 -1960 -2369 1960
rect -6369 -2000 -2369 -1960
rect -2050 1960 1950 2000
rect -2050 -1960 -2010 1960
rect 1910 -1960 1950 1960
rect -2050 -2000 1950 -1960
rect 2269 1960 6269 2000
rect 2269 -1960 2309 1960
rect 6229 -1960 6269 1960
rect 2269 -2000 6269 -1960
rect -6369 -2340 -2369 -2300
rect -6369 -6260 -6329 -2340
rect -2409 -6260 -2369 -2340
rect -6369 -6300 -2369 -6260
rect -2050 -2340 1950 -2300
rect -2050 -6260 -2010 -2340
rect 1910 -6260 1950 -2340
rect -2050 -6300 1950 -6260
rect 2269 -2340 6269 -2300
rect 2269 -6260 2309 -2340
rect 6229 -6260 6269 -2340
rect 2269 -6300 6269 -6260
<< mimcapcontact >>
rect -6329 2340 -2409 6260
rect -2010 2340 1910 6260
rect 2309 2340 6229 6260
rect -6329 -1960 -2409 1960
rect -2010 -1960 1910 1960
rect 2309 -1960 6229 1960
rect -6329 -6260 -2409 -2340
rect -2010 -6260 1910 -2340
rect 2309 -6260 6229 -2340
<< metal4 >>
rect -4421 6261 -4317 6450
rect -102 6261 2 6450
rect 4217 6261 4321 6450
rect 6337 6388 6441 6450
rect 6337 6372 6464 6388
rect -6330 6260 -2408 6261
rect -6330 2340 -6329 6260
rect -2409 2340 -2408 6260
rect -6330 2339 -2408 2340
rect -2011 6260 1911 6261
rect -2011 2340 -2010 6260
rect 1910 2340 1911 6260
rect -2011 2339 1911 2340
rect 2308 6260 6230 6261
rect 2308 2340 2309 6260
rect 6229 2340 6230 6260
rect 2308 2339 6230 2340
rect -4421 1961 -4317 2339
rect -102 1961 2 2339
rect 4217 1961 4321 2339
rect 6337 2228 6384 6372
rect 6448 2228 6464 6372
rect 6337 2212 6464 2228
rect 6337 2088 6441 2212
rect 6337 2072 6464 2088
rect -6330 1960 -2408 1961
rect -6330 -1960 -6329 1960
rect -2409 -1960 -2408 1960
rect -6330 -1961 -2408 -1960
rect -2011 1960 1911 1961
rect -2011 -1960 -2010 1960
rect 1910 -1960 1911 1960
rect -2011 -1961 1911 -1960
rect 2308 1960 6230 1961
rect 2308 -1960 2309 1960
rect 6229 -1960 6230 1960
rect 2308 -1961 6230 -1960
rect -4421 -2339 -4317 -1961
rect -102 -2339 2 -1961
rect 4217 -2339 4321 -1961
rect 6337 -2072 6384 2072
rect 6448 -2072 6464 2072
rect 6337 -2088 6464 -2072
rect 6337 -2212 6441 -2088
rect 6337 -2228 6464 -2212
rect -6330 -2340 -2408 -2339
rect -6330 -6260 -6329 -2340
rect -2409 -6260 -2408 -2340
rect -6330 -6261 -2408 -6260
rect -2011 -2340 1911 -2339
rect -2011 -6260 -2010 -2340
rect 1910 -6260 1911 -2340
rect -2011 -6261 1911 -6260
rect 2308 -2340 6230 -2339
rect 2308 -6260 2309 -2340
rect 6229 -6260 6230 -2340
rect 2308 -6261 6230 -6260
rect -4421 -6450 -4317 -6261
rect -102 -6450 2 -6261
rect 4217 -6450 4321 -6261
rect 6337 -6372 6384 -2228
rect 6448 -6372 6464 -2228
rect 6337 -6388 6464 -6372
rect 6337 -6450 6441 -6388
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 2169 2200 6369 6400
string parameters w 20 l 20 val 815.2 carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
