* NGSPICE file created from top_pll_v1.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_1_MACBVW VSUBS m3_n2650_n13200# m3_n7969_n2600# m3_7988_8000#
+ m3_2669_n7900# m3_n13288_n2600# m3_n2650_2700# m3_2669_2700# m3_n13288_n13200# m3_n7969_n13200#
+ m3_n13288_8000# m3_7988_2700# m3_n2650_n7900# m3_7988_n7900# m3_2669_n13200# m3_n7969_8000#
+ m3_n13288_2700# m3_n7969_n7900# m3_n13288_n7900# m3_2669_n2600# m3_n7969_2700# m3_7988_n13200#
+ c1_n13188_n13100# m3_7988_n2600# m3_n2650_n2600# m3_n2650_8000# m3_2669_8000#
X0 c1_n13188_n13100# m3_2669_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X1 c1_n13188_n13100# m3_n2650_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X2 c1_n13188_n13100# m3_2669_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X3 c1_n13188_n13100# m3_n13288_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X4 c1_n13188_n13100# m3_n7969_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X5 c1_n13188_n13100# m3_n13288_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X6 c1_n13188_n13100# m3_2669_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X7 c1_n13188_n13100# m3_7988_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X8 c1_n13188_n13100# m3_2669_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X9 c1_n13188_n13100# m3_7988_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X10 c1_n13188_n13100# m3_n7969_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X11 c1_n13188_n13100# m3_7988_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X12 c1_n13188_n13100# m3_n7969_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X13 c1_n13188_n13100# m3_7988_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X14 c1_n13188_n13100# m3_n13288_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X15 c1_n13188_n13100# m3_n7969_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X16 c1_n13188_n13100# m3_n2650_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X17 c1_n13188_n13100# m3_n2650_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X18 c1_n13188_n13100# m3_n2650_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X19 c1_n13188_n13100# m3_7988_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X20 c1_n13188_n13100# m3_n13288_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X21 c1_n13188_n13100# m3_n13288_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X22 c1_n13188_n13100# m3_n7969_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X23 c1_n13188_n13100# m3_n2650_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X24 c1_n13188_n13100# m3_2669_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
C0 m3_n2650_n13200# c1_n13188_n13100# 58.61fF
C1 m3_n13288_8000# m3_n7969_8000# 2.73fF
C2 m3_7988_2700# m3_7988_8000# 3.39fF
C3 m3_2669_n2600# m3_n2650_n2600# 2.73fF
C4 m3_n7969_n7900# c1_n13188_n13100# 58.86fF
C5 m3_7988_n7900# m3_2669_n7900# 2.73fF
C6 c1_n13188_n13100# m3_n7969_n2600# 58.86fF
C7 c1_n13188_n13100# m3_7988_n2600# 61.01fF
C8 m3_2669_8000# m3_n2650_8000# 2.73fF
C9 m3_n7969_2700# m3_n7969_n2600# 3.28fF
C10 m3_n2650_n7900# m3_2669_n7900# 2.73fF
C11 m3_2669_n2600# m3_2669_2700# 3.28fF
C12 m3_7988_n2600# m3_7988_2700# 3.39fF
C13 c1_n13188_n13100# m3_n2650_2700# 58.86fF
C14 c1_n13188_n13100# m3_n13288_n2600# 58.61fF
C15 m3_7988_n2600# m3_7988_n7900# 3.39fF
C16 m3_n7969_2700# m3_n2650_2700# 2.73fF
C17 m3_n2650_n13200# m3_n2650_n7900# 3.28fF
C18 c1_n13188_n13100# m3_n7969_8000# 58.61fF
C19 m3_n13288_8000# c1_n13188_n13100# 58.36fF
C20 m3_n7969_n7900# m3_n2650_n7900# 2.73fF
C21 m3_2669_n2600# m3_2669_n7900# 3.28fF
C22 m3_n7969_2700# m3_n7969_8000# 3.28fF
C23 c1_n13188_n13100# m3_n7969_n13200# 58.61fF
C24 c1_n13188_n13100# m3_2669_n13200# 58.61fF
C25 m3_2669_n2600# m3_7988_n2600# 2.73fF
C26 m3_n7969_n13200# m3_n13288_n13200# 2.73fF
C27 m3_n2650_2700# m3_n2650_8000# 3.28fF
C28 m3_n7969_2700# c1_n13188_n13100# 58.86fF
C29 m3_2669_2700# m3_2669_8000# 3.28fF
C30 m3_n2650_8000# m3_n7969_8000# 2.73fF
C31 c1_n13188_n13100# m3_7988_2700# 61.01fF
C32 c1_n13188_n13100# m3_7988_n7900# 61.01fF
C33 c1_n13188_n13100# m3_n13288_n13200# 58.36fF
C34 m3_n13288_n2600# m3_n13288_2700# 3.28fF
C35 m3_2669_8000# m3_7988_8000# 2.73fF
C36 m3_7988_n13200# m3_2669_n13200# 2.73fF
C37 m3_n2650_n2600# m3_n7969_n2600# 2.73fF
C38 m3_n13288_8000# m3_n13288_2700# 3.28fF
C39 c1_n13188_n13100# m3_n2650_n7900# 58.86fF
C40 m3_7988_n13200# c1_n13188_n13100# 60.75fF
C41 m3_n7969_n7900# m3_n13288_n7900# 2.73fF
C42 m3_n2650_2700# m3_n2650_n2600# 3.28fF
C43 c1_n13188_n13100# m3_n2650_8000# 58.61fF
C44 m3_2669_n2600# c1_n13188_n13100# 58.86fF
C45 m3_7988_n13200# m3_7988_n7900# 3.39fF
C46 c1_n13188_n13100# m3_n13288_2700# 58.61fF
C47 m3_n2650_2700# m3_2669_2700# 2.73fF
C48 m3_n13288_n2600# m3_n13288_n7900# 3.28fF
C49 m3_n7969_2700# m3_n13288_2700# 2.73fF
C50 m3_n7969_n7900# m3_n7969_n2600# 3.28fF
C51 c1_n13188_n13100# m3_n2650_n2600# 58.86fF
C52 c1_n13188_n13100# m3_2669_8000# 58.61fF
C53 m3_n13288_n2600# m3_n7969_n2600# 2.73fF
C54 c1_n13188_n13100# m3_n13288_n7900# 58.61fF
C55 c1_n13188_n13100# m3_2669_2700# 58.86fF
C56 m3_2669_n13200# m3_2669_n7900# 3.28fF
C57 m3_n2650_n13200# m3_n7969_n13200# 2.73fF
C58 m3_n7969_n7900# m3_n7969_n13200# 3.28fF
C59 m3_n2650_n7900# m3_n2650_n2600# 3.28fF
C60 c1_n13188_n13100# m3_2669_n7900# 58.86fF
C61 m3_2669_2700# m3_7988_2700# 2.73fF
C62 c1_n13188_n13100# m3_7988_8000# 60.75fF
C63 m3_n2650_n13200# m3_2669_n13200# 2.73fF
C64 m3_n13288_n7900# m3_n13288_n13200# 3.28fF
C65 c1_n13188_n13100# VSUBS 2.51fF
C66 m3_7988_n13200# VSUBS 12.57fF
C67 m3_2669_n13200# VSUBS 12.37fF
C68 m3_n2650_n13200# VSUBS 12.37fF
C69 m3_n7969_n13200# VSUBS 12.37fF
C70 m3_n13288_n13200# VSUBS 12.37fF
C71 m3_7988_n7900# VSUBS 12.57fF
C72 m3_2669_n7900# VSUBS 12.37fF
C73 m3_n2650_n7900# VSUBS 12.37fF
C74 m3_n7969_n7900# VSUBS 12.37fF
C75 m3_n13288_n7900# VSUBS 12.37fF
C76 m3_7988_n2600# VSUBS 12.57fF
C77 m3_2669_n2600# VSUBS 12.37fF
C78 m3_n2650_n2600# VSUBS 12.37fF
C79 m3_n7969_n2600# VSUBS 12.37fF
C80 m3_n13288_n2600# VSUBS 12.37fF
C81 m3_7988_2700# VSUBS 12.57fF
C82 m3_2669_2700# VSUBS 12.37fF
C83 m3_n2650_2700# VSUBS 12.37fF
C84 m3_n7969_2700# VSUBS 12.37fF
C85 m3_n13288_2700# VSUBS 12.37fF
C86 m3_7988_8000# VSUBS 12.57fF
C87 m3_2669_8000# VSUBS 12.37fF
C88 m3_n2650_8000# VSUBS 12.37fF
C89 m3_n7969_8000# VSUBS 12.37fF
C90 m3_n13288_8000# VSUBS 12.37fF
.ends

.subckt cap1_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_MACBVW_0 VSUBS out out out out out out out out out out
+ out out out out out out out out out out out in out out out out sky130_fd_pr__cap_mim_m3_1_MACBVW
C0 out in 2.17fF
C1 in VSUBS -10.03fF
C2 out VSUBS 62.40fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_W3JTNJ VSUBS m3_n6469_n2100# c1_n6369_n6300# m3_2169_n6400#
+ m3_n2150_n6400# c1_2269_n6300# m3_n6469_2200# m3_n2150_n2100# c1_n2050_n6300# m3_n2150_2200#
+ m3_n6469_n6400#
X0 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2 c1_n2050_n6300# m3_n2150_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 c1_n6369_n6300# m3_n6469_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X4 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X5 c1_n6369_n6300# m3_n6469_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X6 c1_n2050_n6300# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X7 c1_n2050_n6300# m3_n2150_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X8 c1_n6369_n6300# m3_n6469_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
C0 m3_n2150_2200# c1_n2050_n6300# 38.10fF
C1 c1_2269_n6300# m3_2169_n6400# 121.67fF
C2 m3_n6469_2200# m3_n2150_2200# 1.75fF
C3 m3_n2150_n2100# m3_2169_n6400# 1.75fF
C4 m3_n2150_n6400# c1_n2050_n6300# 38.10fF
C5 m3_n6469_n2100# m3_n6469_2200# 2.63fF
C6 m3_n6469_n6400# m3_n2150_n6400# 1.75fF
C7 m3_n6469_n2100# m3_n6469_n6400# 2.63fF
C8 m3_n2150_n2100# m3_n2150_2200# 2.63fF
C9 c1_n6369_n6300# m3_n6469_n2100# 38.10fF
C10 c1_n6369_n6300# c1_n2050_n6300# 1.99fF
C11 c1_2269_n6300# c1_n2050_n6300# 1.99fF
C12 c1_n6369_n6300# m3_n6469_2200# 38.10fF
C13 m3_n2150_2200# m3_2169_n6400# 1.75fF
C14 c1_n6369_n6300# m3_n6469_n6400# 38.10fF
C15 m3_n2150_n2100# m3_n2150_n6400# 2.63fF
C16 m3_n2150_n2100# m3_n6469_n2100# 1.75fF
C17 m3_n2150_n2100# c1_n2050_n6300# 38.10fF
C18 m3_n2150_n6400# m3_2169_n6400# 1.75fF
C19 c1_2269_n6300# VSUBS 0.16fF
C20 c1_n2050_n6300# VSUBS 0.16fF
C21 c1_n6369_n6300# VSUBS 0.16fF
C22 m3_n2150_n6400# VSUBS 8.68fF
C23 m3_n6469_n6400# VSUBS 8.68fF
C24 m3_n2150_n2100# VSUBS 8.68fF
C25 m3_n6469_n2100# VSUBS 8.68fF
C26 m3_2169_n6400# VSUBS 26.86fF
C27 m3_n2150_2200# VSUBS 8.68fF
C28 m3_n6469_2200# VSUBS 8.68fF
.ends

.subckt cap2_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_W3JTNJ_0 VSUBS out in out out in out out in out out sky130_fd_pr__cap_mim_m3_1_W3JTNJ
C0 in out 8.08fF
C1 in VSUBS -16.59fF
C2 out VSUBS 13.00fF
.ends

.subckt sky130_fd_pr__res_high_po_5p73_X44RQA a_n573_2292# w_n739_n2890# a_n573_n2724#
X0 a_n573_n2724# a_n573_2292# w_n739_n2890# sky130_fd_pr__res_high_po_5p73 l=2.292e+07u
C0 a_n573_n2724# w_n739_n2890# 1.98fF
C1 a_n573_2292# w_n739_n2890# 1.98fF
.ends

.subckt res_loop_filter vss out in
Xsky130_fd_pr__res_high_po_5p73_X44RQA_0 in vss out sky130_fd_pr__res_high_po_5p73_X44RQA
C0 out vss 3.87fF
C1 in vss 3.02fF
.ends

.subckt loop_filter vc_pex in vss
Xcap1_loop_filter_0 vss vc_pex vss cap1_loop_filter
Xcap2_loop_filter_0 vss in vss cap2_loop_filter
Xres_loop_filter_0 vss res_loop_filter_2/out in res_loop_filter
Xres_loop_filter_1 vss res_loop_filter_2/out vc_pex res_loop_filter
Xres_loop_filter_2 vss res_loop_filter_2/out vc_pex res_loop_filter
C0 in vc_pex 0.18fF
C1 vc_pex vss -38.13fF
C2 res_loop_filter_2/out vss 8.49fF
C3 in vss -18.79fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4ML9WA VSUBS a_429_n486# w_n2457_n634# a_887_n486#
+ a_n29_n486# a_1345_n486# a_n2261_n512# a_1803_n486# a_n487_n486# a_n945_n486# a_n2319_n486#
+ a_n1403_n486# a_2261_n486# a_n1861_n486#
X0 a_2261_n486# a_n2261_n512# a_1803_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X1 a_n945_n486# a_n2261_n512# a_n1403_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X2 a_429_n486# a_n2261_n512# a_n29_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X3 a_1803_n486# a_n2261_n512# a_1345_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X4 a_887_n486# a_n2261_n512# a_429_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X5 a_n487_n486# a_n2261_n512# a_n945_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X6 a_n1403_n486# a_n2261_n512# a_n1861_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X7 a_n1861_n486# a_n2261_n512# a_n2319_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X8 a_n29_n486# a_n2261_n512# a_n487_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X9 a_1345_n486# a_n2261_n512# a_887_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
C0 w_n2457_n634# a_1803_n486# 0.02fF
C1 w_n2457_n634# a_2261_n486# 0.02fF
C2 a_n945_n486# w_n2457_n634# 0.02fF
C3 w_n2457_n634# a_n1861_n486# 0.02fF
C4 w_n2457_n634# a_1345_n486# 0.02fF
C5 w_n2457_n634# a_429_n486# 0.02fF
C6 a_n2319_n486# w_n2457_n634# 0.02fF
C7 w_n2457_n634# a_n1403_n486# 0.02fF
C8 w_n2457_n634# a_n29_n486# 0.02fF
C9 w_n2457_n634# a_n487_n486# 0.02fF
C10 w_n2457_n634# a_887_n486# 0.02fF
C11 a_2261_n486# VSUBS 0.03fF
C12 a_1803_n486# VSUBS 0.03fF
C13 a_1345_n486# VSUBS 0.03fF
C14 a_887_n486# VSUBS 0.03fF
C15 a_429_n486# VSUBS 0.03fF
C16 a_n29_n486# VSUBS 0.03fF
C17 a_n487_n486# VSUBS 0.03fF
C18 a_n945_n486# VSUBS 0.03fF
C19 a_n1403_n486# VSUBS 0.03fF
C20 a_n1861_n486# VSUBS 0.03fF
C21 a_n2319_n486# VSUBS 0.03fF
C22 a_n2261_n512# VSUBS 4.27fF
C23 w_n2457_n634# VSUBS 21.34fF
.ends

.subckt sky130_fd_pr__nfet_01v8_YCGG98 a_n1041_n75# a_n561_n75# a_1167_n75# a_303_n75#
+ a_687_n75# a_n849_n75# a_n369_n75# a_975_n75# a_111_n75# a_495_n75# a_n1137_n75#
+ a_n657_n75# a_n177_n75# a_783_n75# a_n945_n75# a_n465_n75# a_207_n75# a_1071_n75#
+ a_591_n75# a_15_n75# a_n753_n75# w_n1367_n285# a_n273_n75# a_879_n75# a_399_n75#
+ a_n1229_n75# a_n81_n75# a_n1167_n101#
X0 a_207_n75# a_n1167_n101# a_111_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_303_n75# a_n1167_n101# a_207_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_399_n75# a_n1167_n101# a_303_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_495_n75# a_n1167_n101# a_399_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_591_n75# a_n1167_n101# a_495_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_783_n75# a_n1167_n101# a_687_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_687_n75# a_n1167_n101# a_591_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_879_n75# a_n1167_n101# a_783_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_975_n75# a_n1167_n101# a_879_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_n1041_n75# a_n1167_n101# a_n1137_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_n1137_n75# a_n1167_n101# a_n1229_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n561_n75# a_n1167_n101# a_n657_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_1071_n75# a_n1167_n101# a_975_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n945_n75# a_n1167_n101# a_n1041_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n753_n75# a_n1167_n101# a_n849_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n657_n75# a_n1167_n101# a_n753_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n465_n75# a_n1167_n101# a_n561_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n369_n75# a_n1167_n101# a_n465_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_1167_n75# a_n1167_n101# a_1071_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n849_n75# a_n1167_n101# a_n945_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X20 a_15_n75# a_n1167_n101# a_n81_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X21 a_n81_n75# a_n1167_n101# a_n177_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X22 a_111_n75# a_n1167_n101# a_15_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X23 a_n273_n75# a_n1167_n101# a_n369_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X24 a_n177_n75# a_n1167_n101# a_n273_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
C0 a_n1041_n75# a_n657_n75# 0.03fF
C1 a_687_n75# a_591_n75# 0.22fF
C2 a_15_n75# a_111_n75# 0.22fF
C3 a_n945_n75# a_n1137_n75# 0.08fF
C4 a_n753_n75# a_n657_n75# 0.22fF
C5 a_687_n75# a_879_n75# 0.08fF
C6 a_687_n75# a_399_n75# 0.05fF
C7 a_879_n75# a_1071_n75# 0.08fF
C8 a_n465_n75# a_n273_n75# 0.08fF
C9 a_303_n75# a_495_n75# 0.08fF
C10 a_n561_n75# a_n177_n75# 0.03fF
C11 a_n81_n75# a_303_n75# 0.03fF
C12 a_1167_n75# a_879_n75# 0.05fF
C13 a_975_n75# a_591_n75# 0.03fF
C14 a_783_n75# a_687_n75# 0.22fF
C15 a_207_n75# a_591_n75# 0.03fF
C16 a_975_n75# a_879_n75# 0.22fF
C17 a_783_n75# a_1071_n75# 0.05fF
C18 a_n945_n75# a_n657_n75# 0.05fF
C19 a_207_n75# a_399_n75# 0.08fF
C20 a_687_n75# a_495_n75# 0.08fF
C21 a_n1229_n75# a_n849_n75# 0.03fF
C22 a_n465_n75# a_n849_n75# 0.03fF
C23 a_n81_n75# a_n369_n75# 0.05fF
C24 a_783_n75# a_1167_n75# 0.03fF
C25 a_783_n75# a_975_n75# 0.08fF
C26 a_n1041_n75# a_n849_n75# 0.08fF
C27 a_n177_n75# a_n369_n75# 0.08fF
C28 a_n753_n75# a_n849_n75# 0.22fF
C29 a_n1041_n75# a_n1229_n75# 0.08fF
C30 a_207_n75# a_495_n75# 0.05fF
C31 a_111_n75# a_399_n75# 0.05fF
C32 a_15_n75# a_399_n75# 0.03fF
C33 a_n81_n75# a_207_n75# 0.05fF
C34 a_n753_n75# a_n465_n75# 0.05fF
C35 a_207_n75# a_n177_n75# 0.03fF
C36 a_n753_n75# a_n1041_n75# 0.05fF
C37 a_n561_n75# a_n369_n75# 0.08fF
C38 a_n81_n75# a_n273_n75# 0.08fF
C39 a_n945_n75# a_n849_n75# 0.22fF
C40 a_495_n75# a_111_n75# 0.03fF
C41 a_n81_n75# a_111_n75# 0.08fF
C42 a_n657_n75# a_n561_n75# 0.22fF
C43 a_n1229_n75# a_n945_n75# 0.05fF
C44 a_n273_n75# a_n177_n75# 0.22fF
C45 a_n81_n75# a_15_n75# 0.22fF
C46 a_303_n75# a_687_n75# 0.03fF
C47 a_111_n75# a_n177_n75# 0.05fF
C48 a_15_n75# a_n177_n75# 0.08fF
C49 a_n1041_n75# a_n945_n75# 0.22fF
C50 a_879_n75# a_591_n75# 0.05fF
C51 a_399_n75# a_591_n75# 0.08fF
C52 a_n753_n75# a_n945_n75# 0.08fF
C53 a_n81_n75# a_n465_n75# 0.03fF
C54 a_687_n75# a_1071_n75# 0.03fF
C55 a_303_n75# a_207_n75# 0.22fF
C56 a_n273_n75# a_n561_n75# 0.05fF
C57 a_n465_n75# a_n177_n75# 0.05fF
C58 a_n657_n75# a_n369_n75# 0.05fF
C59 a_783_n75# a_591_n75# 0.08fF
C60 a_1167_n75# a_1071_n75# 0.22fF
C61 a_783_n75# a_879_n75# 0.22fF
C62 a_975_n75# a_687_n75# 0.05fF
C63 a_783_n75# a_399_n75# 0.03fF
C64 a_975_n75# a_1071_n75# 0.22fF
C65 a_495_n75# a_591_n75# 0.22fF
C66 a_495_n75# a_879_n75# 0.03fF
C67 a_n849_n75# a_n561_n75# 0.05fF
C68 a_495_n75# a_399_n75# 0.22fF
C69 a_303_n75# a_111_n75# 0.08fF
C70 a_15_n75# a_303_n75# 0.05fF
C71 a_1167_n75# a_975_n75# 0.08fF
C72 a_n465_n75# a_n561_n75# 0.22fF
C73 a_n273_n75# a_n369_n75# 0.22fF
C74 a_783_n75# a_495_n75# 0.05fF
C75 a_n849_n75# a_n1137_n75# 0.05fF
C76 a_n273_n75# a_n657_n75# 0.03fF
C77 a_15_n75# a_n369_n75# 0.03fF
C78 a_n1229_n75# a_n1137_n75# 0.22fF
C79 a_n753_n75# a_n561_n75# 0.08fF
C80 a_n1041_n75# a_n1137_n75# 0.22fF
C81 a_n465_n75# a_n369_n75# 0.22fF
C82 a_207_n75# a_111_n75# 0.22fF
C83 a_15_n75# a_207_n75# 0.08fF
C84 a_n657_n75# a_n849_n75# 0.08fF
C85 a_n753_n75# a_n1137_n75# 0.03fF
C86 a_n81_n75# a_n177_n75# 0.22fF
C87 a_303_n75# a_591_n75# 0.05fF
C88 a_n465_n75# a_n657_n75# 0.08fF
C89 a_n945_n75# a_n561_n75# 0.03fF
C90 a_303_n75# a_399_n75# 0.22fF
C91 a_n273_n75# a_111_n75# 0.03fF
C92 a_n753_n75# a_n369_n75# 0.03fF
C93 a_15_n75# a_n273_n75# 0.05fF
C94 a_1167_n75# w_n1367_n285# 0.10fF
C95 a_1071_n75# w_n1367_n285# 0.07fF
C96 a_975_n75# w_n1367_n285# 0.06fF
C97 a_879_n75# w_n1367_n285# 0.05fF
C98 a_783_n75# w_n1367_n285# 0.04fF
C99 a_687_n75# w_n1367_n285# 0.04fF
C100 a_591_n75# w_n1367_n285# 0.04fF
C101 a_495_n75# w_n1367_n285# 0.04fF
C102 a_399_n75# w_n1367_n285# 0.04fF
C103 a_303_n75# w_n1367_n285# 0.04fF
C104 a_207_n75# w_n1367_n285# 0.04fF
C105 a_111_n75# w_n1367_n285# 0.04fF
C106 a_15_n75# w_n1367_n285# 0.04fF
C107 a_n81_n75# w_n1367_n285# 0.04fF
C108 a_n177_n75# w_n1367_n285# 0.04fF
C109 a_n273_n75# w_n1367_n285# 0.04fF
C110 a_n369_n75# w_n1367_n285# 0.04fF
C111 a_n465_n75# w_n1367_n285# 0.04fF
C112 a_n561_n75# w_n1367_n285# 0.04fF
C113 a_n657_n75# w_n1367_n285# 0.04fF
C114 a_n753_n75# w_n1367_n285# 0.04fF
C115 a_n849_n75# w_n1367_n285# 0.04fF
C116 a_n945_n75# w_n1367_n285# 0.04fF
C117 a_n1041_n75# w_n1367_n285# 0.04fF
C118 a_n1137_n75# w_n1367_n285# 0.04fF
C119 a_n1229_n75# w_n1367_n285# 0.04fF
C120 a_n1167_n101# w_n1367_n285# 2.55fF
.ends

.subckt sky130_fd_pr__nfet_01v8_MUHGM9 a_33_n101# a_n129_n75# a_735_n75# a_255_n75#
+ a_n417_n75# a_n989_n75# a_63_n75# a_543_n75# a_n705_n75# a_n225_n75# a_n33_n75#
+ a_831_n75# a_351_n75# a_n927_n101# a_n513_n75# a_n897_n75# w_n1127_n285# a_639_n75#
+ a_159_n75# a_n801_n75# a_n321_n75# a_927_n75# a_447_n75# a_n609_n75#
X0 a_63_n75# a_33_n101# a_n33_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_927_n75# a_33_n101# a_831_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_n33_n75# a_n927_n101# a_n129_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_159_n75# a_33_n101# a_63_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_255_n75# a_33_n101# a_159_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_351_n75# a_33_n101# a_255_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_447_n75# a_33_n101# a_351_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_543_n75# a_33_n101# a_447_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_735_n75# a_33_n101# a_639_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_831_n75# a_33_n101# a_735_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_639_n75# a_33_n101# a_543_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n321_n75# a_n927_n101# a_n417_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_n801_n75# a_n927_n101# a_n897_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n705_n75# a_n927_n101# a_n801_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n513_n75# a_n927_n101# a_n609_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n417_n75# a_n927_n101# a_n513_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n225_n75# a_n927_n101# a_n321_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n129_n75# a_n927_n101# a_n225_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_n897_n75# a_n927_n101# a_n989_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n609_n75# a_n927_n101# a_n705_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
C0 a_n513_n75# a_n417_n75# 0.22fF
C1 a_255_n75# a_351_n75# 0.22fF
C2 a_735_n75# a_927_n75# 0.08fF
C3 a_159_n75# a_447_n75# 0.05fF
C4 a_351_n75# a_63_n75# 0.05fF
C5 a_543_n75# a_735_n75# 0.08fF
C6 a_n225_n75# a_n33_n75# 0.08fF
C7 a_447_n75# a_831_n75# 0.03fF
C8 a_159_n75# a_n225_n75# 0.03fF
C9 a_n321_n75# a_63_n75# 0.03fF
C10 a_33_n101# a_n927_n101# 0.08fF
C11 a_n321_n75# a_n129_n75# 0.08fF
C12 a_543_n75# a_927_n75# 0.03fF
C13 a_351_n75# a_n33_n75# 0.03fF
C14 a_159_n75# a_351_n75# 0.08fF
C15 a_831_n75# a_639_n75# 0.08fF
C16 a_n321_n75# a_n33_n75# 0.05fF
C17 a_n417_n75# a_n129_n75# 0.05fF
C18 a_n513_n75# a_n129_n75# 0.03fF
C19 a_255_n75# a_543_n75# 0.05fF
C20 a_447_n75# a_639_n75# 0.08fF
C21 a_n33_n75# a_n417_n75# 0.03fF
C22 a_351_n75# a_447_n75# 0.22fF
C23 a_735_n75# a_831_n75# 0.22fF
C24 a_n801_n75# a_n609_n75# 0.08fF
C25 a_255_n75# a_63_n75# 0.08fF
C26 a_n225_n75# a_n609_n75# 0.03fF
C27 a_n801_n75# a_n989_n75# 0.08fF
C28 a_255_n75# a_n129_n75# 0.03fF
C29 a_n897_n75# a_n801_n75# 0.22fF
C30 a_n129_n75# a_63_n75# 0.08fF
C31 a_159_n75# a_543_n75# 0.03fF
C32 a_n609_n75# a_n989_n75# 0.03fF
C33 a_927_n75# a_831_n75# 0.22fF
C34 a_n801_n75# a_n705_n75# 0.22fF
C35 a_n225_n75# a_n321_n75# 0.22fF
C36 a_735_n75# a_447_n75# 0.05fF
C37 a_543_n75# a_831_n75# 0.05fF
C38 a_351_n75# a_639_n75# 0.05fF
C39 a_255_n75# a_n33_n75# 0.05fF
C40 a_n897_n75# a_n609_n75# 0.05fF
C41 a_n897_n75# a_n989_n75# 0.22fF
C42 a_159_n75# a_255_n75# 0.22fF
C43 a_n609_n75# a_n321_n75# 0.05fF
C44 a_n609_n75# a_n705_n75# 0.22fF
C45 a_n33_n75# a_63_n75# 0.22fF
C46 a_n705_n75# a_n989_n75# 0.05fF
C47 a_159_n75# a_63_n75# 0.22fF
C48 a_n801_n75# a_n417_n75# 0.03fF
C49 a_n33_n75# a_n129_n75# 0.22fF
C50 a_n225_n75# a_n417_n75# 0.08fF
C51 a_n513_n75# a_n801_n75# 0.05fF
C52 a_n513_n75# a_n225_n75# 0.05fF
C53 a_159_n75# a_n129_n75# 0.05fF
C54 a_n897_n75# a_n705_n75# 0.08fF
C55 a_543_n75# a_447_n75# 0.22fF
C56 a_735_n75# a_639_n75# 0.22fF
C57 a_n321_n75# a_n705_n75# 0.03fF
C58 a_n609_n75# a_n417_n75# 0.08fF
C59 a_735_n75# a_351_n75# 0.03fF
C60 a_n513_n75# a_n609_n75# 0.22fF
C61 a_255_n75# a_447_n75# 0.08fF
C62 a_159_n75# a_n33_n75# 0.08fF
C63 a_927_n75# a_639_n75# 0.05fF
C64 a_447_n75# a_63_n75# 0.03fF
C65 a_n897_n75# a_n513_n75# 0.03fF
C66 a_543_n75# a_639_n75# 0.22fF
C67 a_n321_n75# a_n417_n75# 0.22fF
C68 a_n417_n75# a_n705_n75# 0.05fF
C69 a_n513_n75# a_n705_n75# 0.08fF
C70 a_n513_n75# a_n321_n75# 0.08fF
C71 a_n225_n75# a_63_n75# 0.05fF
C72 a_543_n75# a_351_n75# 0.08fF
C73 a_n225_n75# a_n129_n75# 0.22fF
C74 a_255_n75# a_639_n75# 0.03fF
C75 a_927_n75# w_n1127_n285# 0.04fF
C76 a_831_n75# w_n1127_n285# 0.04fF
C77 a_735_n75# w_n1127_n285# 0.04fF
C78 a_639_n75# w_n1127_n285# 0.04fF
C79 a_543_n75# w_n1127_n285# 0.04fF
C80 a_447_n75# w_n1127_n285# 0.04fF
C81 a_351_n75# w_n1127_n285# 0.04fF
C82 a_255_n75# w_n1127_n285# 0.04fF
C83 a_159_n75# w_n1127_n285# 0.04fF
C84 a_63_n75# w_n1127_n285# 0.04fF
C85 a_n33_n75# w_n1127_n285# 0.04fF
C86 a_n129_n75# w_n1127_n285# 0.04fF
C87 a_n225_n75# w_n1127_n285# 0.04fF
C88 a_n321_n75# w_n1127_n285# 0.04fF
C89 a_n417_n75# w_n1127_n285# 0.04fF
C90 a_n513_n75# w_n1127_n285# 0.04fF
C91 a_n609_n75# w_n1127_n285# 0.04fF
C92 a_n705_n75# w_n1127_n285# 0.04fF
C93 a_n801_n75# w_n1127_n285# 0.04fF
C94 a_n897_n75# w_n1127_n285# 0.04fF
C95 a_n989_n75# w_n1127_n285# 0.04fF
C96 a_33_n101# w_n1127_n285# 0.99fF
C97 a_n927_n101# w_n1127_n285# 0.99fF
.ends

.subckt sky130_fd_pr__pfet_01v8_NKZXKB VSUBS a_33_n247# a_n801_n150# a_n417_n150#
+ a_351_n150# a_255_n150# a_n705_n150# a_n609_n150# a_159_n150# a_543_n150# a_447_n150#
+ a_831_n150# a_n897_n150# a_n33_n150# a_735_n150# a_n927_n247# a_639_n150# a_n321_n150#
+ a_927_n150# a_n225_n150# a_63_n150# a_n989_n150# a_n513_n150# a_n129_n150# w_n1127_n369#
X0 a_n513_n150# a_n927_n247# a_n609_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_63_n150# a_33_n247# a_n33_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_735_n150# a_33_n247# a_639_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n801_n150# a_n927_n247# a_n897_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n927_n247# a_n225_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n927_n247# a_n513_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_639_n150# a_33_n247# a_543_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n705_n150# a_n927_n247# a_n801_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n33_n150# a_n927_n247# a_n129_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_351_n150# a_33_n247# a_255_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_n609_n150# a_n927_n247# a_n705_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n897_n150# a_n927_n247# a_n989_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_927_n150# a_33_n247# a_831_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_255_n150# a_33_n247# a_159_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n321_n150# a_n927_n247# a_n417_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_543_n150# a_33_n247# a_447_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_831_n150# a_33_n247# a_735_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_159_n150# a_33_n247# a_63_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_n225_n150# a_n927_n247# a_n321_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_447_n150# a_33_n247# a_351_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_159_n150# a_63_n150# 0.43fF
C1 a_n129_n150# a_63_n150# 0.16fF
C2 a_n801_n150# a_n989_n150# 0.16fF
C3 a_255_n150# a_351_n150# 0.43fF
C4 a_n513_n150# a_n417_n150# 0.43fF
C5 a_n609_n150# a_n321_n150# 0.10fF
C6 a_927_n150# a_543_n150# 0.07fF
C7 a_n225_n150# a_n33_n150# 0.16fF
C8 a_543_n150# a_735_n150# 0.16fF
C9 a_n321_n150# a_n705_n150# 0.07fF
C10 a_n609_n150# a_n989_n150# 0.07fF
C11 a_447_n150# a_63_n150# 0.07fF
C12 a_n801_n150# a_n417_n150# 0.07fF
C13 a_447_n150# a_639_n150# 0.16fF
C14 a_831_n150# a_639_n150# 0.16fF
C15 a_n989_n150# a_n705_n150# 0.10fF
C16 a_n33_n150# a_63_n150# 0.43fF
C17 a_927_n150# a_831_n150# 0.43fF
C18 a_n609_n150# a_n417_n150# 0.16fF
C19 a_351_n150# a_63_n150# 0.10fF
C20 a_255_n150# a_63_n150# 0.16fF
C21 a_735_n150# a_831_n150# 0.43fF
C22 a_447_n150# a_735_n150# 0.10fF
C23 a_351_n150# a_639_n150# 0.10fF
C24 a_255_n150# a_639_n150# 0.07fF
C25 a_n417_n150# a_n705_n150# 0.10fF
C26 a_n513_n150# a_n225_n150# 0.10fF
C27 a_n225_n150# a_63_n150# 0.10fF
C28 a_n513_n150# a_n897_n150# 0.07fF
C29 a_n321_n150# a_n129_n150# 0.16fF
C30 a_735_n150# a_351_n150# 0.07fF
C31 a_n417_n150# a_n321_n150# 0.43fF
C32 a_543_n150# a_159_n150# 0.07fF
C33 a_n897_n150# a_n801_n150# 0.43fF
C34 a_n513_n150# a_n801_n150# 0.10fF
C35 a_n609_n150# a_n225_n150# 0.07fF
C36 a_159_n150# a_n129_n150# 0.10fF
C37 a_543_n150# a_447_n150# 0.43fF
C38 a_543_n150# a_831_n150# 0.10fF
C39 a_n33_n150# a_n321_n150# 0.10fF
C40 a_n609_n150# a_n897_n150# 0.10fF
C41 a_n417_n150# a_n129_n150# 0.10fF
C42 a_n609_n150# a_n513_n150# 0.43fF
C43 a_927_n150# a_639_n150# 0.10fF
C44 a_159_n150# a_447_n150# 0.10fF
C45 a_n897_n150# a_n705_n150# 0.16fF
C46 a_n513_n150# a_n705_n150# 0.16fF
C47 a_735_n150# a_639_n150# 0.43fF
C48 a_543_n150# a_351_n150# 0.16fF
C49 a_255_n150# a_543_n150# 0.10fF
C50 a_n225_n150# a_n321_n150# 0.43fF
C51 a_n33_n150# a_159_n150# 0.16fF
C52 a_n33_n150# a_n129_n150# 0.43fF
C53 a_n609_n150# a_n801_n150# 0.16fF
C54 a_447_n150# a_831_n150# 0.07fF
C55 a_927_n150# a_735_n150# 0.16fF
C56 a_159_n150# a_351_n150# 0.16fF
C57 a_n33_n150# a_n417_n150# 0.07fF
C58 a_255_n150# a_159_n150# 0.43fF
C59 a_255_n150# a_n129_n150# 0.07fF
C60 a_n801_n150# a_n705_n150# 0.43fF
C61 a_33_n247# a_n927_n247# 0.09fF
C62 a_n513_n150# a_n321_n150# 0.16fF
C63 a_n321_n150# a_63_n150# 0.07fF
C64 a_n897_n150# a_n989_n150# 0.43fF
C65 a_n225_n150# a_159_n150# 0.07fF
C66 a_n225_n150# a_n129_n150# 0.43fF
C67 a_447_n150# a_351_n150# 0.43fF
C68 a_255_n150# a_447_n150# 0.16fF
C69 a_n609_n150# a_n705_n150# 0.43fF
C70 a_n225_n150# a_n417_n150# 0.16fF
C71 a_543_n150# a_639_n150# 0.43fF
C72 a_n33_n150# a_351_n150# 0.07fF
C73 a_n513_n150# a_n129_n150# 0.07fF
C74 a_255_n150# a_n33_n150# 0.10fF
C75 a_927_n150# VSUBS 0.03fF
C76 a_831_n150# VSUBS 0.03fF
C77 a_735_n150# VSUBS 0.03fF
C78 a_639_n150# VSUBS 0.03fF
C79 a_543_n150# VSUBS 0.03fF
C80 a_447_n150# VSUBS 0.03fF
C81 a_351_n150# VSUBS 0.03fF
C82 a_255_n150# VSUBS 0.03fF
C83 a_159_n150# VSUBS 0.03fF
C84 a_63_n150# VSUBS 0.03fF
C85 a_n33_n150# VSUBS 0.03fF
C86 a_n129_n150# VSUBS 0.03fF
C87 a_n225_n150# VSUBS 0.03fF
C88 a_n321_n150# VSUBS 0.03fF
C89 a_n417_n150# VSUBS 0.03fF
C90 a_n513_n150# VSUBS 0.03fF
C91 a_n609_n150# VSUBS 0.03fF
C92 a_n705_n150# VSUBS 0.03fF
C93 a_n801_n150# VSUBS 0.03fF
C94 a_n897_n150# VSUBS 0.03fF
C95 a_n989_n150# VSUBS 0.03fF
C96 a_33_n247# VSUBS 1.04fF
C97 a_n927_n247# VSUBS 1.04fF
C98 w_n1127_n369# VSUBS 6.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_8GRULZ a_n1761_n132# a_1045_n44# a_n1461_n44# a_n1103_n44#
+ a_n29_n44# a_n387_n44# a_1761_n44# a_n1819_n44# a_1403_n44# a_687_n44# w_n1957_n254#
+ a_329_n44# a_n745_n44#
X0 a_329_n44# a_n1761_n132# a_n29_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X1 a_1761_n44# a_n1761_n132# a_1403_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X2 a_n745_n44# a_n1761_n132# a_n1103_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X3 a_1045_n44# a_n1761_n132# a_687_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X4 a_n29_n44# a_n1761_n132# a_n387_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X5 a_n1103_n44# a_n1761_n132# a_n1461_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X6 a_n387_n44# a_n1761_n132# a_n745_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X7 a_687_n44# a_n1761_n132# a_329_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X8 a_1403_n44# a_n1761_n132# a_1045_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X9 a_n1461_n44# a_n1761_n132# a_n1819_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
C0 a_687_n44# a_329_n44# 0.04fF
C1 a_1045_n44# a_1403_n44# 0.04fF
C2 a_n387_n44# a_n29_n44# 0.04fF
C3 a_n1461_n44# a_n1819_n44# 0.04fF
C4 a_n745_n44# a_n387_n44# 0.04fF
C5 a_n745_n44# a_n1103_n44# 0.04fF
C6 a_n1461_n44# a_n1103_n44# 0.04fF
C7 a_n29_n44# a_329_n44# 0.04fF
C8 a_1045_n44# a_687_n44# 0.04fF
C9 a_1761_n44# a_1403_n44# 0.04fF
C10 a_1761_n44# w_n1957_n254# 0.04fF
C11 a_1403_n44# w_n1957_n254# 0.04fF
C12 a_1045_n44# w_n1957_n254# 0.04fF
C13 a_687_n44# w_n1957_n254# 0.04fF
C14 a_329_n44# w_n1957_n254# 0.04fF
C15 a_n29_n44# w_n1957_n254# 0.04fF
C16 a_n387_n44# w_n1957_n254# 0.04fF
C17 a_n745_n44# w_n1957_n254# 0.04fF
C18 a_n1103_n44# w_n1957_n254# 0.04fF
C19 a_n1461_n44# w_n1957_n254# 0.04fF
C20 a_n1819_n44# w_n1957_n254# 0.04fF
C21 a_n1761_n132# w_n1957_n254# 3.23fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ND88ZC VSUBS a_303_n150# a_n753_n150# a_n369_n150#
+ w_n1367_n369# a_207_n150# a_n657_n150# a_591_n150# a_n1229_n150# a_n945_n150# a_495_n150#
+ a_n1041_n150# a_n849_n150# a_n81_n150# a_399_n150# a_783_n150# a_1071_n150# a_687_n150#
+ a_975_n150# a_n1137_n150# a_n273_n150# a_111_n150# a_879_n150# a_n177_n150# a_n561_n150#
+ a_15_n150# a_1167_n150# a_n1167_n247# a_n465_n150#
X0 a_n1137_n150# a_n1167_n247# a_n1229_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_495_n150# a_n1167_n247# a_399_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n561_n150# a_n1167_n247# a_n657_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_111_n150# a_n1167_n247# a_15_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_783_n150# a_n1167_n247# a_687_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_1071_n150# a_n1167_n247# a_975_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_399_n150# a_n1167_n247# a_303_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n465_n150# a_n1167_n247# a_n561_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_687_n150# a_n1167_n247# a_591_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n753_n150# a_n1167_n247# a_n849_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_975_n150# a_n1167_n247# a_879_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n81_n150# a_n1167_n247# a_n177_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_15_n150# a_n1167_n247# a_n81_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_n1041_n150# a_n1167_n247# a_n1137_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n369_n150# a_n1167_n247# a_n465_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_n657_n150# a_n1167_n247# a_n753_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_879_n150# a_n1167_n247# a_783_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_n945_n150# a_n1167_n247# a_n1041_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_1167_n150# a_n1167_n247# a_1071_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_303_n150# a_n1167_n247# a_207_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X20 a_n273_n150# a_n1167_n247# a_n369_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X21 a_591_n150# a_n1167_n247# a_495_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X22 a_n849_n150# a_n1167_n247# a_n945_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_207_n150# a_n1167_n247# a_111_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X24 a_n177_n150# a_n1167_n247# a_n273_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_399_n150# a_783_n150# 0.07fF
C1 a_15_n150# a_n369_n150# 0.07fF
C2 a_n561_n150# a_n465_n150# 0.43fF
C3 a_n81_n150# a_303_n150# 0.07fF
C4 a_879_n150# a_687_n150# 0.16fF
C5 a_n657_n150# a_n369_n150# 0.10fF
C6 w_n1367_n369# a_975_n150# 0.05fF
C7 a_111_n150# a_207_n150# 0.43fF
C8 a_591_n150# a_783_n150# 0.16fF
C9 a_975_n150# a_1167_n150# 0.16fF
C10 a_879_n150# a_495_n150# 0.07fF
C11 a_399_n150# a_207_n150# 0.16fF
C12 a_n369_n150# a_n753_n150# 0.07fF
C13 a_n81_n150# a_n177_n150# 0.43fF
C14 a_303_n150# a_15_n150# 0.10fF
C15 a_n657_n150# a_n1041_n150# 0.07fF
C16 a_879_n150# w_n1367_n369# 0.04fF
C17 a_1071_n150# a_975_n150# 0.43fF
C18 a_879_n150# a_1167_n150# 0.10fF
C19 a_591_n150# a_207_n150# 0.07fF
C20 a_783_n150# a_975_n150# 0.16fF
C21 a_n81_n150# a_n465_n150# 0.07fF
C22 a_n1137_n150# a_n945_n150# 0.16fF
C23 a_n1041_n150# a_n753_n150# 0.10fF
C24 a_n561_n150# a_n849_n150# 0.10fF
C25 a_15_n150# a_n177_n150# 0.16fF
C26 a_399_n150# a_111_n150# 0.10fF
C27 a_n273_n150# a_111_n150# 0.07fF
C28 a_879_n150# a_1071_n150# 0.16fF
C29 a_879_n150# a_783_n150# 0.43fF
C30 a_n849_n150# a_n945_n150# 0.43fF
C31 a_n657_n150# a_n465_n150# 0.16fF
C32 a_591_n150# a_399_n150# 0.16fF
C33 a_n1229_n150# a_n945_n150# 0.10fF
C34 a_n81_n150# a_207_n150# 0.10fF
C35 a_n465_n150# a_n753_n150# 0.10fF
C36 a_n561_n150# a_n273_n150# 0.10fF
C37 a_n1137_n150# a_n753_n150# 0.07fF
C38 a_687_n150# a_495_n150# 0.16fF
C39 a_303_n150# a_687_n150# 0.07fF
C40 a_207_n150# a_15_n150# 0.16fF
C41 a_n369_n150# a_n177_n150# 0.16fF
C42 a_n657_n150# a_n849_n150# 0.16fF
C43 a_303_n150# a_495_n150# 0.16fF
C44 a_n81_n150# a_111_n150# 0.16fF
C45 a_n465_n150# a_n369_n150# 0.43fF
C46 a_591_n150# a_975_n150# 0.07fF
C47 a_n849_n150# a_n753_n150# 0.43fF
C48 a_n273_n150# a_n81_n150# 0.16fF
C49 a_111_n150# a_15_n150# 0.43fF
C50 a_n561_n150# a_n945_n150# 0.07fF
C51 a_399_n150# a_15_n150# 0.07fF
C52 a_n273_n150# a_15_n150# 0.10fF
C53 a_879_n150# a_591_n150# 0.10fF
C54 a_n657_n150# a_n273_n150# 0.07fF
C55 a_1071_n150# a_687_n150# 0.07fF
C56 w_n1367_n369# a_1167_n150# 0.14fF
C57 a_687_n150# a_783_n150# 0.43fF
C58 a_n1041_n150# a_n1137_n150# 0.43fF
C59 a_783_n150# a_495_n150# 0.10fF
C60 a_n465_n150# a_n177_n150# 0.10fF
C61 a_879_n150# a_975_n150# 0.43fF
C62 a_n657_n150# a_n561_n150# 0.43fF
C63 a_1071_n150# w_n1367_n369# 0.07fF
C64 a_n1041_n150# a_n849_n150# 0.16fF
C65 a_1071_n150# a_1167_n150# 0.43fF
C66 a_783_n150# a_1167_n150# 0.07fF
C67 a_207_n150# a_495_n150# 0.10fF
C68 a_303_n150# a_207_n150# 0.43fF
C69 a_n561_n150# a_n753_n150# 0.16fF
C70 a_n1041_n150# a_n1229_n150# 0.16fF
C71 a_n657_n150# a_n945_n150# 0.10fF
C72 a_n273_n150# a_n369_n150# 0.43fF
C73 a_n81_n150# a_15_n150# 0.43fF
C74 a_1071_n150# a_783_n150# 0.10fF
C75 a_207_n150# a_n177_n150# 0.07fF
C76 a_n753_n150# a_n945_n150# 0.16fF
C77 a_111_n150# a_495_n150# 0.07fF
C78 a_303_n150# a_111_n150# 0.16fF
C79 a_n849_n150# a_n465_n150# 0.07fF
C80 a_399_n150# a_687_n150# 0.10fF
C81 a_399_n150# a_495_n150# 0.43fF
C82 a_399_n150# a_303_n150# 0.43fF
C83 a_n561_n150# a_n369_n150# 0.16fF
C84 a_n849_n150# a_n1137_n150# 0.10fF
C85 a_111_n150# a_n177_n150# 0.10fF
C86 a_591_n150# a_687_n150# 0.43fF
C87 a_591_n150# a_495_n150# 0.43fF
C88 a_591_n150# a_303_n150# 0.10fF
C89 a_n273_n150# a_n177_n150# 0.43fF
C90 a_n1137_n150# a_n1229_n150# 0.43fF
C91 a_n657_n150# a_n753_n150# 0.43fF
C92 a_n273_n150# a_n465_n150# 0.16fF
C93 a_n81_n150# a_n369_n150# 0.10fF
C94 a_687_n150# a_975_n150# 0.10fF
C95 a_n1041_n150# a_n945_n150# 0.43fF
C96 a_n849_n150# a_n1229_n150# 0.07fF
C97 a_n561_n150# a_n177_n150# 0.07fF
C98 a_1167_n150# VSUBS 0.03fF
C99 a_1071_n150# VSUBS 0.03fF
C100 a_975_n150# VSUBS 0.03fF
C101 a_879_n150# VSUBS 0.03fF
C102 a_783_n150# VSUBS 0.03fF
C103 a_687_n150# VSUBS 0.03fF
C104 a_591_n150# VSUBS 0.03fF
C105 a_495_n150# VSUBS 0.03fF
C106 a_399_n150# VSUBS 0.03fF
C107 a_303_n150# VSUBS 0.03fF
C108 a_207_n150# VSUBS 0.03fF
C109 a_111_n150# VSUBS 0.03fF
C110 a_15_n150# VSUBS 0.03fF
C111 a_n81_n150# VSUBS 0.03fF
C112 a_n177_n150# VSUBS 0.03fF
C113 a_n273_n150# VSUBS 0.03fF
C114 a_n369_n150# VSUBS 0.03fF
C115 a_n465_n150# VSUBS 0.03fF
C116 a_n561_n150# VSUBS 0.03fF
C117 a_n657_n150# VSUBS 0.03fF
C118 a_n753_n150# VSUBS 0.03fF
C119 a_n849_n150# VSUBS 0.03fF
C120 a_n945_n150# VSUBS 0.03fF
C121 a_n1041_n150# VSUBS 0.03fF
C122 a_n1137_n150# VSUBS 0.03fF
C123 a_n1229_n150# VSUBS 0.03fF
C124 a_n1167_n247# VSUBS 2.63fF
C125 w_n1367_n369# VSUBS 7.85fF
.ends

.subckt charge_pump nswitch vdd nUp vss Down biasp out pswitch iref nDown Up
Xsky130_fd_pr__pfet_01v8_4ML9WA_0 vss pswitch vdd pswitch pswitch pswitch nUp pswitch
+ pswitch pswitch pswitch pswitch pswitch pswitch sky130_fd_pr__pfet_01v8_4ML9WA
Xsky130_fd_pr__nfet_01v8_YCGG98_0 vss out out vss vss vss out out vss vss out vss
+ out out out vss out vss out out out vss vss vss out vss vss nswitch sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_1 iref vss vss iref iref iref vss vss iref iref vss
+ iref vss vss vss iref vss iref vss vss vss vss iref iref vss iref iref iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_2 biasp vss vss biasp biasp biasp vss vss biasp biasp
+ vss biasp vss vss vss biasp vss biasp vss vss vss vss biasp biasp vss biasp biasp
+ iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_MUHGM9_0 nDown iref nswitch vss nswitch nswitch vss nswitch
+ iref nswitch nswitch vss nswitch Down iref iref vss vss nswitch nswitch iref nswitch
+ vss nswitch sky130_fd_pr__nfet_01v8_MUHGM9
Xsky130_fd_pr__pfet_01v8_NKZXKB_0 vss Up pswitch pswitch pswitch vdd biasp pswitch
+ pswitch pswitch vdd vdd biasp pswitch pswitch nUp vdd biasp pswitch pswitch vdd
+ pswitch biasp biasp vdd sky130_fd_pr__pfet_01v8_NKZXKB
Xsky130_fd_pr__nfet_01v8_8GRULZ_0 Down nswitch nswitch nswitch nswitch nswitch nswitch
+ nswitch nswitch nswitch vss nswitch nswitch sky130_fd_pr__nfet_01v8_8GRULZ
Xsky130_fd_pr__pfet_01v8_ND88ZC_0 vss vdd out out vdd out vdd out vdd out vdd vdd
+ vdd vdd out out vdd vdd out out vdd vdd vdd out out out out pswitch vdd sky130_fd_pr__pfet_01v8_ND88ZC
Xsky130_fd_pr__pfet_01v8_ND88ZC_1 vss biasp vdd vdd vdd vdd biasp vdd biasp vdd biasp
+ biasp biasp biasp vdd vdd biasp biasp vdd vdd biasp biasp biasp vdd vdd vdd vdd
+ biasp biasp sky130_fd_pr__pfet_01v8_ND88ZC
C0 nswitch out 1.28fF
C1 nswitch Down 2.27fF
C2 biasp pswitch 3.11fF
C3 vdd pswitch 3.98fF
C4 nDown Down 0.13fF
C5 nDown nswitch 0.31fF
C6 nswitch iref 1.91fF
C7 Up pswitch 0.70fF
C8 vdd out 6.66fF
C9 nUp Up 0.15fF
C10 biasp nswitch 0.03fF
C11 nswitch vdd 0.07fF
C12 nUp pswitch 5.66fF
C13 biasp iref 0.80fF
C14 pswitch out 4.91fF
C15 nUp out 0.31fF
C16 nswitch pswitch 0.06fF
C17 biasp vdd 2.64fF
C18 nUp Down 0.25fF
C19 vdd vss 35.71fF
C20 Down vss 4.77fF
C21 Up vss 1.17fF
C22 nswitch vss 6.39fF
C23 nDown vss 1.11fF
C24 biasp vss 8.73fF
C25 iref vss 10.12fF
C26 out vss -3.49fF
C27 pswitch vss 3.45fF
C28 nUp vss 5.85fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4798MH VSUBS a_81_n156# a_111_n125# a_15_n125# a_n173_n125#
+ w_n311_n344# a_n111_n156# a_n15_n156# a_n81_n125#
X0 a_n81_n125# a_n111_n156# a_n173_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n15_n156# a_n81_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_81_n156# a_15_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n173_n125# a_111_n125# 0.08fF
C1 a_15_n125# a_111_n125# 0.36fF
C2 w_n311_n344# a_n81_n125# 0.09fF
C3 a_15_n125# a_n173_n125# 0.13fF
C4 a_n81_n125# a_111_n125# 0.13fF
C5 a_n81_n125# a_n173_n125# 0.36fF
C6 a_15_n125# a_n81_n125# 0.36fF
C7 w_n311_n344# a_111_n125# 0.14fF
C8 w_n311_n344# a_n173_n125# 0.14fF
C9 a_15_n125# w_n311_n344# 0.09fF
C10 a_81_n156# a_n15_n156# 0.02fF
C11 a_n111_n156# a_n15_n156# 0.02fF
C12 a_111_n125# VSUBS 0.03fF
C13 a_15_n125# VSUBS 0.03fF
C14 a_n81_n125# VSUBS 0.03fF
C15 a_n173_n125# VSUBS 0.03fF
C16 a_81_n156# VSUBS 0.05fF
C17 a_n15_n156# VSUBS 0.05fF
C18 a_n111_n156# VSUBS 0.05fF
C19 w_n311_n344# VSUBS 2.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_BHR94T a_n15_n151# w_n311_n335# a_81_n151# a_111_n125#
+ a_15_n125# a_n173_n125# a_n111_n151# a_n81_n125#
X0 a_111_n125# a_81_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n15_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n15_n151# a_n111_n151# 0.02fF
C1 a_n81_n125# a_111_n125# 0.13fF
C2 a_n173_n125# a_111_n125# 0.08fF
C3 a_15_n125# a_111_n125# 0.36fF
C4 a_81_n151# a_n15_n151# 0.02fF
C5 a_n173_n125# a_n81_n125# 0.36fF
C6 a_15_n125# a_n81_n125# 0.36fF
C7 a_n173_n125# a_15_n125# 0.13fF
C8 a_111_n125# w_n311_n335# 0.17fF
C9 a_15_n125# w_n311_n335# 0.12fF
C10 a_n81_n125# w_n311_n335# 0.12fF
C11 a_n173_n125# w_n311_n335# 0.17fF
C12 a_81_n151# w_n311_n335# 0.05fF
C13 a_n15_n151# w_n311_n335# 0.05fF
C14 a_n111_n151# w_n311_n335# 0.05fF
.ends

.subckt trans_gate m1_187_n605# m1_45_n513# vss vdd
Xsky130_fd_pr__pfet_01v8_4798MH_0 vss vss m1_187_n605# m1_45_n513# m1_45_n513# vdd
+ vss vss m1_187_n605# sky130_fd_pr__pfet_01v8_4798MH
Xsky130_fd_pr__nfet_01v8_BHR94T_0 vdd vss vdd m1_187_n605# m1_45_n513# m1_45_n513#
+ vdd m1_187_n605# sky130_fd_pr__nfet_01v8_BHR94T
C0 vdd m1_187_n605# 0.55fF
C1 m1_187_n605# m1_45_n513# 0.36fF
C2 vdd m1_45_n513# 0.69fF
C3 m1_187_n605# vss 0.93fF
C4 m1_45_n513# vss 1.31fF
C5 vdd vss 3.36fF
.ends

.subckt sky130_fd_pr__pfet_01v8_7KT7MH VSUBS a_n111_n186# a_111_n125# a_15_n125# a_n173_n125#
+ w_n311_n344# a_n81_n125#
X0 a_n81_n125# a_n111_n186# a_n173_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n111_n186# a_n81_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_n111_n186# a_15_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_111_n125# w_n311_n344# 0.14fF
C1 a_n81_n125# w_n311_n344# 0.09fF
C2 a_15_n125# w_n311_n344# 0.09fF
C3 a_111_n125# a_n81_n125# 0.13fF
C4 w_n311_n344# a_n173_n125# 0.14fF
C5 a_111_n125# a_15_n125# 0.36fF
C6 a_n81_n125# a_15_n125# 0.36fF
C7 a_111_n125# a_n173_n125# 0.08fF
C8 a_n81_n125# a_n173_n125# 0.36fF
C9 a_15_n125# a_n173_n125# 0.13fF
C10 a_111_n125# VSUBS 0.03fF
C11 a_15_n125# VSUBS 0.03fF
C12 a_n81_n125# VSUBS 0.03fF
C13 a_n173_n125# VSUBS 0.03fF
C14 a_n111_n186# VSUBS 0.26fF
C15 w_n311_n344# VSUBS 2.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS6QM w_n311_n335# a_111_n125# a_15_n125# a_n173_n125#
+ a_n111_n151# a_n81_n125#
X0 a_111_n125# a_n111_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n111_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_15_n125# a_n173_n125# 0.13fF
C1 a_15_n125# a_111_n125# 0.36fF
C2 a_111_n125# a_n173_n125# 0.08fF
C3 a_15_n125# a_n81_n125# 0.36fF
C4 a_n173_n125# a_n81_n125# 0.36fF
C5 a_111_n125# a_n81_n125# 0.13fF
C6 a_111_n125# w_n311_n335# 0.17fF
C7 a_15_n125# w_n311_n335# 0.12fF
C8 a_n81_n125# w_n311_n335# 0.12fF
C9 a_n173_n125# w_n311_n335# 0.17fF
C10 a_n111_n151# w_n311_n335# 0.25fF
.ends

.subckt inverter_cp_x1 out in vss vdd
Xsky130_fd_pr__pfet_01v8_7KT7MH_0 vss in out vdd vdd vdd out sky130_fd_pr__pfet_01v8_7KT7MH
Xsky130_fd_pr__nfet_01v8_2BS6QM_0 vss out vss vss in out sky130_fd_pr__nfet_01v8_2BS6QM
C0 out vdd 0.10fF
C1 out in 0.32fF
C2 out vss 0.77fF
C3 in vss 0.95fF
C4 vdd vss 3.13fF
.ends

.subckt clock_inverter vss inverter_cp_x1_2/in CLK vdd inverter_cp_x1_0/out CLK_d
+ nCLK_d
Xtrans_gate_0 nCLK_d inverter_cp_x1_0/out vss vdd trans_gate
Xinverter_cp_x1_0 inverter_cp_x1_0/out CLK vss vdd inverter_cp_x1
Xinverter_cp_x1_1 inverter_cp_x1_2/in CLK vss vdd inverter_cp_x1
Xinverter_cp_x1_2 CLK_d inverter_cp_x1_2/in vss vdd inverter_cp_x1
C0 inverter_cp_x1_2/in CLK 0.31fF
C1 vdd CLK_d 0.03fF
C2 vdd inverter_cp_x1_0/out 0.28fF
C3 vdd CLK 0.36fF
C4 vdd inverter_cp_x1_2/in 0.21fF
C5 nCLK_d inverter_cp_x1_0/out 0.11fF
C6 vdd nCLK_d 0.03fF
C7 CLK_d inverter_cp_x1_2/in 0.12fF
C8 CLK inverter_cp_x1_0/out 0.31fF
C9 CLK_d vss 0.96fF
C10 inverter_cp_x1_2/in vss 2.01fF
C11 inverter_cp_x1_0/out vss 1.97fF
C12 CLK vss 3.03fF
C13 nCLK_d vss 1.44fF
C14 vdd vss 16.51fF
.ends

.subckt sky130_fd_pr__pfet_01v8_MJG8BZ VSUBS a_n125_n95# a_63_n95# w_n263_n314# a_n33_n95#
+ a_n63_n192#
X0 a_63_n95# a_n63_n192# a_n33_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n33_n95# a_n63_n192# a_n125_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
C0 a_63_n95# a_n125_n95# 0.10fF
C1 a_63_n95# a_n33_n95# 0.28fF
C2 a_n125_n95# a_n33_n95# 0.28fF
C3 w_n263_n314# a_63_n95# 0.11fF
C4 w_n263_n314# a_n125_n95# 0.11fF
C5 w_n263_n314# a_n33_n95# 0.08fF
C6 a_63_n95# VSUBS 0.03fF
C7 a_n33_n95# VSUBS 0.03fF
C8 a_n125_n95# VSUBS 0.03fF
C9 a_n63_n192# VSUBS 0.20fF
C10 w_n263_n314# VSUBS 1.80fF
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS854 w_n311_n335# a_n129_n213# a_111_n125# a_15_n125#
+ a_n173_n125# a_n81_n125#
X0 a_111_n125# a_n129_n213# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n129_n213# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n129_n213# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n81_n125# a_n173_n125# 0.36fF
C1 a_111_n125# a_n81_n125# 0.13fF
C2 a_15_n125# a_n173_n125# 0.13fF
C3 a_111_n125# a_15_n125# 0.36fF
C4 a_n81_n125# a_15_n125# 0.36fF
C5 a_n129_n213# a_n173_n125# 0.02fF
C6 a_n129_n213# a_111_n125# 0.01fF
C7 a_n129_n213# a_n81_n125# 0.10fF
C8 a_n129_n213# a_15_n125# 0.10fF
C9 a_111_n125# a_n173_n125# 0.08fF
C10 a_111_n125# w_n311_n335# 0.05fF
C11 a_15_n125# w_n311_n335# 0.05fF
C12 a_n81_n125# w_n311_n335# 0.05fF
C13 a_n173_n125# w_n311_n335# 0.05fF
C14 a_n129_n213# w_n311_n335# 0.49fF
.ends

.subckt sky130_fd_pr__nfet_01v8_KU9PSX a_n125_n95# a_n33_n95# a_n81_n183# w_n263_n305#
X0 a_n33_n95# a_n81_n183# a_n125_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n125_n95# a_n81_n183# a_n33_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
C0 a_n33_n95# a_n125_n95# 0.88fF
C1 a_n81_n183# a_n125_n95# 0.16fF
C2 a_n81_n183# a_n33_n95# 0.10fF
C3 a_n33_n95# w_n263_n305# 0.07fF
C4 a_n125_n95# w_n263_n305# 0.13fF
C5 a_n81_n183# w_n263_n305# 0.31fF
.ends

.subckt latch_diff m1_657_280# nQ Q vss CLK vdd nD D
Xsky130_fd_pr__pfet_01v8_MJG8BZ_0 vss vdd vdd vdd nQ Q sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__pfet_01v8_MJG8BZ_1 vss vdd vdd vdd Q nQ sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__nfet_01v8_2BS854_0 vss CLK vss m1_657_280# m1_657_280# vss sky130_fd_pr__nfet_01v8_2BS854
Xsky130_fd_pr__nfet_01v8_KU9PSX_0 m1_657_280# Q nD vss sky130_fd_pr__nfet_01v8_KU9PSX
Xsky130_fd_pr__nfet_01v8_KU9PSX_1 m1_657_280# nQ D vss sky130_fd_pr__nfet_01v8_KU9PSX
C0 nQ vdd 0.16fF
C1 m1_657_280# Q 0.94fF
C2 m1_657_280# CLK 0.24fF
C3 nD Q 0.05fF
C4 m1_657_280# nQ 1.41fF
C5 D Q 0.05fF
C6 nQ nD 0.05fF
C7 nQ D 0.05fF
C8 nQ Q 0.93fF
C9 vdd Q 0.16fF
C10 nQ vss 1.16fF
C11 D vss 0.53fF
C12 Q vss -0.55fF
C13 m1_657_280# vss 1.88fF
C14 nD vss 0.16fF
C15 CLK vss 0.87fF
C16 vdd vss 5.98fF
.ends

.subckt DFlipFlop latch_diff_0/m1_657_280# vss latch_diff_1/D clock_inverter_0/inverter_cp_x1_2/in
+ nQ Q latch_diff_1/nD D latch_diff_1/m1_657_280# latch_diff_0/D vdd CLK clock_inverter_0/inverter_cp_x1_0/out
+ nCLK latch_diff_0/nD
Xclock_inverter_0 vss clock_inverter_0/inverter_cp_x1_2/in D vdd clock_inverter_0/inverter_cp_x1_0/out
+ latch_diff_0/D latch_diff_0/nD clock_inverter
Xlatch_diff_0 latch_diff_0/m1_657_280# latch_diff_1/nD latch_diff_1/D vss CLK vdd
+ latch_diff_0/nD latch_diff_0/D latch_diff
Xlatch_diff_1 latch_diff_1/m1_657_280# nQ Q vss nCLK vdd latch_diff_1/nD latch_diff_1/D
+ latch_diff
C0 Q latch_diff_1/nD 0.01fF
C1 latch_diff_1/m1_657_280# latch_diff_1/nD 0.42fF
C2 latch_diff_1/m1_657_280# latch_diff_1/D 0.32fF
C3 latch_diff_1/D latch_diff_0/nD 0.41fF
C4 latch_diff_0/D latch_diff_1/nD 0.04fF
C5 latch_diff_0/D latch_diff_1/D 0.11fF
C6 vdd latch_diff_0/nD 0.14fF
C7 latch_diff_1/nD latch_diff_1/D 0.33fF
C8 vdd latch_diff_0/D 0.09fF
C9 latch_diff_1/m1_657_280# latch_diff_0/m1_657_280# 0.18fF
C10 latch_diff_0/m1_657_280# latch_diff_0/nD 0.38fF
C11 latch_diff_0/D latch_diff_0/m1_657_280# 0.37fF
C12 vdd latch_diff_1/nD 0.02fF
C13 vdd latch_diff_1/D 0.03fF
C14 vdd clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C15 nQ latch_diff_1/nD 0.08fF
C16 nQ latch_diff_1/D 0.11fF
C17 latch_diff_0/m1_657_280# latch_diff_1/nD 0.14fF
C18 latch_diff_0/m1_657_280# latch_diff_1/D 0.43fF
C19 nQ vss 0.57fF
C20 Q vss -0.92fF
C21 latch_diff_1/m1_657_280# vss 0.64fF
C22 nCLK vss 0.83fF
C23 latch_diff_1/nD vss 1.83fF
C24 latch_diff_1/D vss -0.30fF
C25 latch_diff_0/m1_657_280# vss 0.72fF
C26 CLK vss 0.83fF
C27 latch_diff_0/D vss 1.29fF
C28 clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C29 clock_inverter_0/inverter_cp_x1_0/out vss 1.84fF
C30 D vss 3.27fF
C31 latch_diff_0/nD vss 1.74fF
C32 vdd vss 32.62fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ZP3U9B VSUBS a_n221_n84# a_159_n84# w_n359_n303# a_n63_n110#
+ a_n129_n84# a_33_n110# a_n159_n110# a_63_n84# a_129_n110# a_n33_n84#
X0 a_n129_n84# a_n159_n110# a_n221_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_63_n84# a_33_n110# a_n33_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_n33_n84# a_n63_n110# a_n129_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_159_n84# a_129_n110# a_63_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_63_n84# a_n33_n84# 0.24fF
C1 w_n359_n303# a_159_n84# 0.08fF
C2 a_n129_n84# a_n221_n84# 0.24fF
C3 a_63_n84# a_159_n84# 0.24fF
C4 a_n33_n84# a_n129_n84# 0.24fF
C5 a_n33_n84# a_n221_n84# 0.09fF
C6 w_n359_n303# a_63_n84# 0.06fF
C7 a_n129_n84# a_159_n84# 0.05fF
C8 a_n221_n84# a_159_n84# 0.04fF
C9 a_n33_n84# a_159_n84# 0.09fF
C10 a_n63_n110# a_n159_n110# 0.02fF
C11 w_n359_n303# a_n129_n84# 0.06fF
C12 w_n359_n303# a_n221_n84# 0.08fF
C13 w_n359_n303# a_n33_n84# 0.05fF
C14 a_33_n110# a_129_n110# 0.02fF
C15 a_63_n84# a_n129_n84# 0.09fF
C16 a_63_n84# a_n221_n84# 0.05fF
C17 a_n63_n110# a_33_n110# 0.02fF
C18 a_159_n84# VSUBS 0.03fF
C19 a_63_n84# VSUBS 0.03fF
C20 a_n33_n84# VSUBS 0.03fF
C21 a_n129_n84# VSUBS 0.03fF
C22 a_n221_n84# VSUBS 0.03fF
C23 a_129_n110# VSUBS 0.05fF
C24 a_33_n110# VSUBS 0.05fF
C25 a_n63_n110# VSUBS 0.05fF
C26 a_n159_n110# VSUBS 0.05fF
C27 w_n359_n303# VSUBS 2.19fF
.ends

.subckt sky130_fd_pr__nfet_01v8_DXA56D w_n359_n252# a_n33_n42# a_129_n68# a_n159_n68#
+ a_n221_n42# a_159_n42# a_n129_n42# a_33_n68# a_n63_n68# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n129_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_159_n42# a_129_n68# a_63_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_n129_n42# a_n159_n68# a_n221_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n129_n42# a_n221_n42# 0.12fF
C1 a_63_n42# a_n33_n42# 0.12fF
C2 a_n221_n42# a_159_n42# 0.02fF
C3 a_n159_n68# a_n63_n68# 0.02fF
C4 a_n129_n42# a_n33_n42# 0.12fF
C5 a_n129_n42# a_63_n42# 0.05fF
C6 a_n33_n42# a_159_n42# 0.05fF
C7 a_63_n42# a_159_n42# 0.12fF
C8 a_33_n68# a_129_n68# 0.02fF
C9 a_n129_n42# a_159_n42# 0.03fF
C10 a_n221_n42# a_n33_n42# 0.05fF
C11 a_n221_n42# a_63_n42# 0.03fF
C12 a_33_n68# a_n63_n68# 0.02fF
C13 a_159_n42# w_n359_n252# 0.07fF
C14 a_63_n42# w_n359_n252# 0.06fF
C15 a_n33_n42# w_n359_n252# 0.06fF
C16 a_n129_n42# w_n359_n252# 0.06fF
C17 a_n221_n42# w_n359_n252# 0.07fF
C18 a_129_n68# w_n359_n252# 0.05fF
C19 a_33_n68# w_n359_n252# 0.05fF
C20 a_n63_n68# w_n359_n252# 0.05fF
C21 a_n159_n68# w_n359_n252# 0.05fF
.ends

.subckt inverter_min_x4 in vss out vdd
Xsky130_fd_pr__pfet_01v8_ZP3U9B_0 vss out out vdd in vdd in in vdd in out sky130_fd_pr__pfet_01v8_ZP3U9B
Xsky130_fd_pr__nfet_01v8_DXA56D_0 vss out in in out out vss in in vss sky130_fd_pr__nfet_01v8_DXA56D
C0 out vdd 0.62fF
C1 out in 0.67fF
C2 in vdd 0.33fF
C3 out vss 0.66fF
C4 in vss 1.89fF
C5 vdd vss 3.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_5RJ8EK a_n33_n42# a_33_n68# w_n263_n252# a_n63_n68#
+ a_n125_n42# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n125_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n33_n42# a_63_n42# 0.12fF
C1 a_n125_n42# a_n33_n42# 0.12fF
C2 a_33_n68# a_n63_n68# 0.02fF
C3 a_n125_n42# a_63_n42# 0.05fF
C4 a_63_n42# w_n263_n252# 0.09fF
C5 a_n33_n42# w_n263_n252# 0.07fF
C6 a_n125_n42# w_n263_n252# 0.09fF
C7 a_33_n68# w_n263_n252# 0.05fF
C8 a_n63_n68# w_n263_n252# 0.05fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ZPB9BB VSUBS a_n63_n110# a_33_n110# a_n125_n84# a_63_n84#
+ w_n263_n303# a_n33_n84#
X0 a_63_n84# a_33_n110# a_n33_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_n33_n84# a_n63_n110# a_n125_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_n63_n110# a_33_n110# 0.02fF
C1 a_n125_n84# a_n33_n84# 0.24fF
C2 w_n263_n303# a_n33_n84# 0.07fF
C3 a_63_n84# a_n125_n84# 0.09fF
C4 a_63_n84# w_n263_n303# 0.10fF
C5 a_63_n84# a_n33_n84# 0.24fF
C6 w_n263_n303# a_n125_n84# 0.10fF
C7 a_63_n84# VSUBS 0.03fF
C8 a_n33_n84# VSUBS 0.03fF
C9 a_n125_n84# VSUBS 0.03fF
C10 a_33_n110# VSUBS 0.05fF
C11 a_n63_n110# VSUBS 0.05fF
C12 w_n263_n303# VSUBS 1.74fF
.ends

.subckt inverter_min_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_5RJ8EK_0 vss in vss in out out sky130_fd_pr__nfet_01v8_5RJ8EK
Xsky130_fd_pr__pfet_01v8_ZPB9BB_0 vss in in out out vdd vdd sky130_fd_pr__pfet_01v8_ZPB9BB
C0 vdd in 0.01fF
C1 vdd out 0.15fF
C2 out in 0.30fF
C3 vdd vss 2.93fF
C4 out vss 0.66fF
C5 in vss 0.72fF
.ends

.subckt div_by_2 vss vdd clock_inverter_0/inverter_cp_x1_2/in CLK_2 nCLK_2 o1 CLK
+ out_div o2 clock_inverter_0/inverter_cp_x1_0/out nout_div
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vss DFlipFlop_0/latch_diff_1/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ nout_div out_div DFlipFlop_0/latch_diff_1/nD nout_div DFlipFlop_0/latch_diff_1/m1_657_280#
+ DFlipFlop_0/latch_diff_0/D vdd DFlipFlop_0/CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_0/nD DFlipFlop
Xclock_inverter_0 vss clock_inverter_0/inverter_cp_x1_2/in CLK vdd clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_0/CLK DFlipFlop_0/nCLK clock_inverter
Xinverter_min_x4_0 o1 vss CLK_2 vdd inverter_min_x4
Xinverter_min_x4_1 o2 vss nCLK_2 vdd inverter_min_x4
Xinverter_min_x2_0 nout_div o2 vss vdd inverter_min_x2
Xinverter_min_x2_1 out_div o1 vss vdd inverter_min_x2
C0 DFlipFlop_0/nCLK vdd 0.30fF
C1 o2 nCLK_2 0.11fF
C2 out_div vdd 0.03fF
C3 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vdd 0.03fF
C4 DFlipFlop_0/latch_diff_1/nD nout_div 1.18fF
C5 DFlipFlop_0/latch_diff_1/m1_657_280# o1 0.02fF
C6 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop_0/CLK 0.29fF
C7 DFlipFlop_0/latch_diff_0/m1_657_280# DFlipFlop_0/CLK 0.26fF
C8 nout_div DFlipFlop_0/latch_diff_0/D 0.09fF
C9 DFlipFlop_0/latch_diff_1/D nout_div 0.64fF
C10 CLK_2 o1 0.11fF
C11 nout_div vdd 0.16fF
C12 o2 vdd 0.14fF
C13 DFlipFlop_0/CLK DFlipFlop_0/latch_diff_0/nD 0.12fF
C14 DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_1/m1_657_280# 0.26fF
C15 nout_div DFlipFlop_0/CLK 0.42fF
C16 DFlipFlop_0/nCLK nout_div 0.43fF
C17 nCLK_2 vdd 0.08fF
C18 nout_div out_div 0.22fF
C19 nout_div DFlipFlop_0/latch_diff_0/m1_657_280# 0.24fF
C20 vdd o1 0.14fF
C21 DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/CLK 0.11fF
C22 DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_1/nD -0.09fF
C23 DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_0/D 0.13fF
C24 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vdd 0.03fF
C25 DFlipFlop_0/latch_diff_1/D DFlipFlop_0/CLK -0.48fF
C26 out_div o1 0.01fF
C27 DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_1/D 0.08fF
C28 DFlipFlop_0/nCLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.46fF
C29 CLK_2 vdd 0.08fF
C30 DFlipFlop_0/latch_diff_1/m1_657_280# nout_div 0.21fF
C31 nout_div DFlipFlop_0/latch_diff_0/nD 0.07fF
C32 DFlipFlop_0/latch_diff_1/m1_657_280# o2 0.02fF
C33 clock_inverter_0/inverter_cp_x1_0/out vdd 0.10fF
C34 DFlipFlop_0/CLK vdd 0.40fF
C35 nCLK_2 vss 1.08fF
C36 o2 vss 2.21fF
C37 CLK_2 vss 1.08fF
C38 o1 vss 2.21fF
C39 DFlipFlop_0/CLK vss 1.03fF
C40 clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C41 clock_inverter_0/inverter_cp_x1_0/out vss 1.85fF
C42 CLK vss 3.27fF
C43 DFlipFlop_0/nCLK vss 1.76fF
C44 out_div vss -0.77fF
C45 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.63fF
C46 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C47 DFlipFlop_0/latch_diff_1/D vss -1.72fF
C48 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C49 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C50 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.89fF
C51 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.80fF
C52 nout_div vss 4.41fF
C53 DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C54 vdd vss 64.43fF
.ends

.subckt sky130_fd_pr__pfet_01v8_58ZKDE VSUBS a_n257_n777# a_n129_n600# a_n221_n600#
+ w_n257_n702#
X0 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X1 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X2 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X3 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
C0 a_n257_n777# a_n221_n600# 0.25fF
C1 a_n257_n777# a_n129_n600# 0.29fF
C2 a_n221_n600# a_n129_n600# 7.87fF
C3 a_n129_n600# VSUBS 0.10fF
C4 a_n221_n600# VSUBS 0.25fF
C5 a_n257_n777# VSUBS 1.05fF
C6 w_n257_n702# VSUBS 2.16fF
.ends

.subckt sky130_fd_pr__nfet_01v8_T69Y3A a_n129_n300# a_n221_n300# w_n257_n327# a_n257_n404#
X0 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
C0 a_n257_n404# a_n221_n300# 0.21fF
C1 a_n221_n300# a_n129_n300# 4.05fF
C2 a_n257_n404# a_n129_n300# 0.30fF
C3 a_n129_n300# w_n257_n327# 0.11fF
C4 a_n221_n300# w_n257_n327# 0.25fF
C5 a_n257_n404# w_n257_n327# 1.11fF
.ends

.subckt buffer_salida a_678_n100# out in vss vdd
Xsky130_fd_pr__pfet_01v8_58ZKDE_1 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_2 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_3 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_0 a_678_n100# vss vss in sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_1 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_4 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_5 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_2 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_3 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_6 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_4 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_7 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_70 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_8 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_5 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_71 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_60 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_6 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_9 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_72 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_61 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_50 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_7 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_62 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_51 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_40 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_8 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_63 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_52 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_41 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_30 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_9 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_20 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_64 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_53 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_42 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_31 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_10 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_21 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_65 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_54 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_43 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_32 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_11 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_22 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_66 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_55 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_44 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_33 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_12 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_23 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_67 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_56 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_45 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_34 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_13 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_24 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_68 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_57 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_46 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_35 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_14 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_69 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_58 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_47 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_36 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_25 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_15 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_59 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_48 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_37 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_26 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_16 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_49 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_38 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_27 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_70 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_17 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_39 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_28 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_71 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_60 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_18 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_29 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_72 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_61 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_50 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_19 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_62 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_51 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_40 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_63 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_52 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_41 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_30 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_20 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_64 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_53 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_42 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_31 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_10 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_21 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_65 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_54 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_43 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_32 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_11 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_22 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_66 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_55 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_44 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_33 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_12 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_23 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_67 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_56 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_45 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_34 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_13 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_24 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_68 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_57 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_46 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_35 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_14 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_69 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_58 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_47 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_36 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_25 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_15 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_59 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_48 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_37 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_26 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_16 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_49 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_38 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_27 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_17 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_39 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_28 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_18 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_29 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_19 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_0 vss in a_678_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
C0 a_3996_n100# vdd 3.68fF
C1 a_678_n100# a_3996_n100# 6.52fF
C2 a_3996_n100# out 55.19fF
C3 a_678_n100# vdd 0.08fF
C4 out vdd 47.17fF
C5 vdd in 0.02fF
C6 a_678_n100# in 0.81fF
C7 vdd vss 20.93fF
C8 out vss 35.17fF
C9 a_3996_n100# vss 49.53fF
C10 a_678_n100# vss 13.08fF
C11 in vss 0.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_CBAU6Y a_n73_n150# a_n33_n238# w_n211_n360# a_15_n150#
X0 a_15_n150# a_n33_n238# a_n73_n150# w_n211_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n33_n238# a_n73_n150# 0.02fF
C1 a_15_n150# a_n33_n238# 0.02fF
C2 a_15_n150# a_n73_n150# 0.51fF
C3 a_15_n150# w_n211_n360# 0.23fF
C4 a_n73_n150# w_n211_n360# 0.23fF
C5 a_n33_n238# w_n211_n360# 0.17fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4757AC VSUBS a_n73_n150# a_n33_181# w_n211_n369# a_15_n150#
X0 a_15_n150# a_n33_181# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n33_181# a_15_n150# 0.01fF
C1 a_n73_n150# a_15_n150# 0.51fF
C2 w_n211_n369# a_n33_181# 0.05fF
C3 a_n73_n150# w_n211_n369# 0.20fF
C4 w_n211_n369# a_15_n150# 0.20fF
C5 a_n73_n150# a_n33_181# 0.01fF
C6 a_15_n150# VSUBS 0.03fF
C7 a_n73_n150# VSUBS 0.03fF
C8 a_n33_181# VSUBS 0.13fF
C9 w_n211_n369# VSUBS 1.98fF
.ends

.subckt sky130_fd_pr__nfet_01v8_7H8F5S a_n465_172# a_n417_n150# a_351_n150# a_255_n150#
+ w_n647_n360# a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150#
X0 a_159_n150# a_n465_172# a_63_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n225_n150# a_n465_172# a_n321_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_447_n150# a_n465_172# a_351_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_63_n150# a_n465_172# a_n33_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n465_172# a_n225_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n465_172# a_n509_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n33_n150# a_n465_172# a_n129_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_351_n150# a_n465_172# a_255_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_255_n150# a_n465_172# a_159_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n321_n150# a_n465_172# a_n417_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n129_n150# a_159_n150# 0.10fF
C1 a_n465_172# a_n129_n150# 0.10fF
C2 a_n509_n150# a_n321_n150# 0.16fF
C3 a_n465_172# a_159_n150# 0.10fF
C4 a_n417_n150# a_n321_n150# 0.43fF
C5 a_63_n150# a_447_n150# 0.07fF
C6 a_63_n150# a_255_n150# 0.16fF
C7 a_n129_n150# a_255_n150# 0.07fF
C8 a_447_n150# a_159_n150# 0.10fF
C9 a_n465_172# a_447_n150# 0.01fF
C10 a_n417_n150# a_n33_n150# 0.07fF
C11 a_255_n150# a_159_n150# 0.43fF
C12 a_n465_172# a_255_n150# 0.10fF
C13 a_351_n150# a_n33_n150# 0.07fF
C14 a_n33_n150# a_n321_n150# 0.10fF
C15 a_447_n150# a_255_n150# 0.16fF
C16 a_n509_n150# a_n225_n150# 0.10fF
C17 a_n129_n150# a_n509_n150# 0.07fF
C18 a_n417_n150# a_n225_n150# 0.16fF
C19 a_n417_n150# a_n129_n150# 0.10fF
C20 a_n465_172# a_n509_n150# 0.01fF
C21 a_351_n150# a_63_n150# 0.10fF
C22 a_n417_n150# a_n465_172# 0.10fF
C23 a_63_n150# a_n321_n150# 0.07fF
C24 a_351_n150# a_159_n150# 0.16fF
C25 a_n225_n150# a_n321_n150# 0.43fF
C26 a_n465_172# a_351_n150# 0.10fF
C27 a_n129_n150# a_n321_n150# 0.16fF
C28 a_n465_172# a_n321_n150# 0.10fF
C29 a_63_n150# a_n33_n150# 0.43fF
C30 a_n33_n150# a_n225_n150# 0.16fF
C31 a_351_n150# a_447_n150# 0.43fF
C32 a_n129_n150# a_n33_n150# 0.43fF
C33 a_351_n150# a_255_n150# 0.43fF
C34 a_n33_n150# a_159_n150# 0.16fF
C35 a_n465_172# a_n33_n150# 0.10fF
C36 a_n33_n150# a_255_n150# 0.10fF
C37 a_63_n150# a_n225_n150# 0.10fF
C38 a_n417_n150# a_n509_n150# 0.43fF
C39 a_n129_n150# a_63_n150# 0.16fF
C40 a_n129_n150# a_n225_n150# 0.43fF
C41 a_63_n150# a_159_n150# 0.43fF
C42 a_n225_n150# a_159_n150# 0.07fF
C43 a_n465_172# a_63_n150# 0.10fF
C44 a_n465_172# a_n225_n150# 0.10fF
C45 a_447_n150# w_n647_n360# 0.17fF
C46 a_351_n150# w_n647_n360# 0.10fF
C47 a_255_n150# w_n647_n360# 0.08fF
C48 a_159_n150# w_n647_n360# 0.07fF
C49 a_63_n150# w_n647_n360# 0.04fF
C50 a_n33_n150# w_n647_n360# 0.04fF
C51 a_n129_n150# w_n647_n360# 0.04fF
C52 a_n225_n150# w_n647_n360# 0.07fF
C53 a_n321_n150# w_n647_n360# 0.08fF
C54 a_n417_n150# w_n647_n360# 0.10fF
C55 a_n509_n150# w_n647_n360# 0.17fF
C56 a_n465_172# w_n647_n360# 1.49fF
.ends

.subckt sky130_fd_pr__pfet_01v8_8DL6ZL VSUBS a_n417_n150# a_351_n150# a_255_n150#
+ a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n465_n247# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150# w_n647_n369#
X0 a_63_n150# a_n465_n247# a_n33_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n129_n150# a_n465_n247# a_n225_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n417_n150# a_n465_n247# a_n509_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n33_n150# a_n465_n247# a_n129_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_351_n150# a_n465_n247# a_255_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_255_n150# a_n465_n247# a_159_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n321_n150# a_n465_n247# a_n417_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_159_n150# a_n465_n247# a_63_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n225_n150# a_n465_n247# a_n321_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_447_n150# a_n465_n247# a_351_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n321_n150# a_n33_n150# 0.10fF
C1 a_n321_n150# a_n129_n150# 0.16fF
C2 a_n321_n150# a_n225_n150# 0.43fF
C3 a_63_n150# a_159_n150# 0.43fF
C4 a_63_n150# a_n33_n150# 0.43fF
C5 a_63_n150# a_n129_n150# 0.16fF
C6 a_n321_n150# w_n647_n369# 0.05fF
C7 a_63_n150# a_n225_n150# 0.10fF
C8 a_63_n150# w_n647_n369# 0.02fF
C9 a_n417_n150# a_n33_n150# 0.07fF
C10 a_n417_n150# a_n129_n150# 0.10fF
C11 a_n465_n247# a_159_n150# 0.08fF
C12 a_n465_n247# a_n33_n150# 0.08fF
C13 a_n417_n150# a_n225_n150# 0.16fF
C14 a_n465_n247# a_n129_n150# 0.08fF
C15 a_n321_n150# a_63_n150# 0.07fF
C16 a_n465_n247# a_n225_n150# 0.08fF
C17 a_n417_n150# w_n647_n369# 0.07fF
C18 a_n465_n247# w_n647_n369# 0.47fF
C19 a_n321_n150# a_n417_n150# 0.43fF
C20 a_255_n150# a_351_n150# 0.43fF
C21 a_n321_n150# a_n465_n247# 0.08fF
C22 a_447_n150# a_255_n150# 0.16fF
C23 a_n465_n247# a_63_n150# 0.08fF
C24 a_n417_n150# a_n465_n247# 0.08fF
C25 a_447_n150# a_351_n150# 0.43fF
C26 a_n509_n150# a_n129_n150# 0.07fF
C27 a_n509_n150# a_n225_n150# 0.10fF
C28 a_255_n150# a_159_n150# 0.43fF
C29 a_255_n150# a_n33_n150# 0.10fF
C30 a_255_n150# a_n129_n150# 0.07fF
C31 a_n509_n150# w_n647_n369# 0.14fF
C32 a_255_n150# w_n647_n369# 0.05fF
C33 a_n321_n150# a_n509_n150# 0.16fF
C34 a_159_n150# a_351_n150# 0.16fF
C35 a_n33_n150# a_351_n150# 0.07fF
C36 a_255_n150# a_63_n150# 0.16fF
C37 a_447_n150# a_159_n150# 0.10fF
C38 a_n509_n150# a_n417_n150# 0.43fF
C39 w_n647_n369# a_351_n150# 0.07fF
C40 a_447_n150# w_n647_n369# 0.14fF
C41 a_255_n150# a_n465_n247# 0.08fF
C42 a_63_n150# a_351_n150# 0.10fF
C43 a_447_n150# a_63_n150# 0.07fF
C44 a_n465_n247# a_351_n150# 0.08fF
C45 a_159_n150# a_n33_n150# 0.16fF
C46 a_n129_n150# a_159_n150# 0.10fF
C47 a_n129_n150# a_n33_n150# 0.43fF
C48 a_159_n150# a_n225_n150# 0.07fF
C49 a_n33_n150# a_n225_n150# 0.16fF
C50 a_n129_n150# a_n225_n150# 0.43fF
C51 a_159_n150# w_n647_n369# 0.04fF
C52 w_n647_n369# a_n33_n150# 0.02fF
C53 a_n129_n150# w_n647_n369# 0.02fF
C54 w_n647_n369# a_n225_n150# 0.04fF
C55 a_447_n150# VSUBS 0.03fF
C56 a_351_n150# VSUBS 0.03fF
C57 a_255_n150# VSUBS 0.03fF
C58 a_159_n150# VSUBS 0.03fF
C59 a_63_n150# VSUBS 0.03fF
C60 a_n33_n150# VSUBS 0.03fF
C61 a_n129_n150# VSUBS 0.03fF
C62 a_n225_n150# VSUBS 0.03fF
C63 a_n321_n150# VSUBS 0.03fF
C64 a_n417_n150# VSUBS 0.03fF
C65 a_n509_n150# VSUBS 0.03fF
C66 a_n465_n247# VSUBS 1.07fF
C67 w_n647_n369# VSUBS 4.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EDT3AT a_15_n11# a_n33_n99# w_n211_n221# a_n73_n11#
X0 a_15_n11# a_n33_n99# a_n73_n11# w_n211_n221# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n33_n99# a_n73_n11# 0.02fF
C1 a_15_n11# a_n73_n11# 0.15fF
C2 a_15_n11# a_n33_n99# 0.02fF
C3 a_15_n11# w_n211_n221# 0.09fF
C4 a_n73_n11# w_n211_n221# 0.09fF
C5 a_n33_n99# w_n211_n221# 0.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AQR2CW a_n33_66# a_n78_n106# w_n216_n254# a_20_n106#
X0 a_20_n106# a_n33_66# a_n78_n106# w_n216_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=200000u
C0 a_20_n106# a_n78_n106# 0.21fF
C1 a_20_n106# w_n216_n254# 0.14fF
C2 a_n78_n106# w_n216_n254# 0.14fF
C3 a_n33_66# w_n216_n254# 0.12fF
.ends

.subckt sky130_fd_pr__pfet_01v8_HRYSXS VSUBS a_n33_n211# a_n78_n114# w_n216_n334#
+ a_20_n114#
X0 a_20_n114# a_n33_n211# a_n78_n114# w_n216_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=200000u
C0 a_n78_n114# a_20_n114# 0.42fF
C1 a_n78_n114# w_n216_n334# 0.20fF
C2 w_n216_n334# a_20_n114# 0.20fF
C3 a_20_n114# VSUBS 0.03fF
C4 a_n78_n114# VSUBS 0.03fF
C5 a_n33_n211# VSUBS 0.12fF
C6 w_n216_n334# VSUBS 1.66fF
.ends

.subckt inverter_csvco in vbulkn out vbulkp vdd vss
Xsky130_fd_pr__nfet_01v8_AQR2CW_0 in vss vbulkn out sky130_fd_pr__nfet_01v8_AQR2CW
Xsky130_fd_pr__pfet_01v8_HRYSXS_0 vbulkn in vdd vbulkp out sky130_fd_pr__pfet_01v8_HRYSXS
C0 in vss 0.01fF
C1 vbulkp vdd 0.04fF
C2 vbulkp out 0.08fF
C3 in vdd 0.01fF
C4 in out 0.11fF
C5 vbulkp vbulkn 2.49fF
C6 out vbulkn 0.60fF
C7 vdd vbulkn 0.06fF
C8 in vbulkn 0.54fF
C9 vss vbulkn 0.17fF
.ends

.subckt csvco_branch vctrl in vbp cap_vco_0/t D0 out inverter_csvco_0/vss vss vdd
+ inverter_csvco_0/vdd
Xsky130_fd_pr__nfet_01v8_7H8F5S_0 vctrl inverter_csvco_0/vss inverter_csvco_0/vss
+ vss vss inverter_csvco_0/vss vss vss inverter_csvco_0/vss vss inverter_csvco_0/vss
+ vss vss sky130_fd_pr__nfet_01v8_7H8F5S
Xsky130_fd_pr__pfet_01v8_8DL6ZL_0 vss inverter_csvco_0/vdd inverter_csvco_0/vdd vdd
+ inverter_csvco_0/vdd vdd vdd inverter_csvco_0/vdd vbp vdd inverter_csvco_0/vdd vdd
+ vdd vdd sky130_fd_pr__pfet_01v8_8DL6ZL
Xsky130_fd_pr__nfet_01v8_EDT3AT_0 cap_vco_0/t D0 vss out sky130_fd_pr__nfet_01v8_EDT3AT
Xinverter_csvco_0 in vss out vdd inverter_csvco_0/vdd inverter_csvco_0/vss inverter_csvco
C0 inverter_csvco_0/vdd out 0.02fF
C1 vbp inverter_csvco_0/vdd 0.75fF
C2 cap_vco_0/t out 0.70fF
C3 inverter_csvco_0/vdd vdd 1.89fF
C4 cap_vco_0/t vdd 0.04fF
C5 inverter_csvco_0/vdd in 0.01fF
C6 D0 out 0.09fF
C7 inverter_csvco_0/vss D0 0.02fF
C8 vbp vdd 1.21fF
C9 out in 0.06fF
C10 vctrl inverter_csvco_0/vss 0.87fF
C11 inverter_csvco_0/vdd cap_vco_0/t 0.10fF
C12 inverter_csvco_0/vss out 0.03fF
C13 inverter_csvco_0/vss in 0.01fF
C14 out vss 0.93fF
C15 inverter_csvco_0/vdd vss 0.26fF
C16 in vss 0.69fF
C17 D0 vss -0.67fF
C18 vbp vss 0.13fF
C19 vdd vss 9.58fF
C20 cap_vco_0/t vss 7.22fF
C21 inverter_csvco_0/vss vss 1.79fF
C22 vctrl vss 3.06fF
.ends

.subckt ring_osc vctrl vdd vss csvco_branch_0/inverter_csvco_0/vss csvco_branch_2/vbp
+ D0 csvco_branch_2/cap_vco_0/t out_vco
Xsky130_fd_pr__nfet_01v8_CBAU6Y_0 vss vctrl vss csvco_branch_2/vbp sky130_fd_pr__nfet_01v8_CBAU6Y
Xsky130_fd_pr__pfet_01v8_4757AC_0 vss vdd csvco_branch_2/vbp vdd csvco_branch_2/vbp
+ sky130_fd_pr__pfet_01v8_4757AC
Xcsvco_branch_0 vctrl out_vco csvco_branch_2/vbp csvco_branch_0/cap_vco_0/t D0 csvco_branch_1/in
+ csvco_branch_0/inverter_csvco_0/vss vss vdd csvco_branch_0/inverter_csvco_0/vdd
+ csvco_branch
Xcsvco_branch_2 vctrl csvco_branch_2/in csvco_branch_2/vbp csvco_branch_2/cap_vco_0/t
+ D0 out_vco csvco_branch_2/inverter_csvco_0/vss vss vdd csvco_branch_2/inverter_csvco_0/vdd
+ csvco_branch
Xcsvco_branch_1 vctrl csvco_branch_1/in csvco_branch_2/vbp csvco_branch_1/cap_vco_0/t
+ D0 csvco_branch_2/in csvco_branch_1/inverter_csvco_0/vss vss vdd csvco_branch_1/inverter_csvco_0/vdd
+ csvco_branch
C0 D0 csvco_branch_2/inverter_csvco_0/vss 0.68fF
C1 csvco_branch_2/in out_vco 0.58fF
C2 csvco_branch_0/inverter_csvco_0/vdd csvco_branch_2/vbp 0.06fF
C3 D0 csvco_branch_1/inverter_csvco_0/vss 0.68fF
C4 csvco_branch_0/inverter_csvco_0/vdd vdd 0.13fF
C5 vdd csvco_branch_1/inverter_csvco_0/vdd 0.19fF
C6 csvco_branch_1/cap_vco_0/t out_vco 0.03fF
C7 vdd csvco_branch_2/inverter_csvco_0/vdd 0.10fF
C8 csvco_branch_0/inverter_csvco_0/vss csvco_branch_2/vbp 0.06fF
C9 out_vco csvco_branch_0/cap_vco_0/t 0.03fF
C10 D0 csvco_branch_0/inverter_csvco_0/vss 0.49fF
C11 csvco_branch_1/in out_vco 0.76fF
C12 vctrl csvco_branch_2/vbp 0.06fF
C13 vdd csvco_branch_2/vbp 1.49fF
C14 D0 vctrl 4.41fF
C15 csvco_branch_2/in vss 1.60fF
C16 csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C17 csvco_branch_1/cap_vco_0/t vss 7.10fF
C18 csvco_branch_1/inverter_csvco_0/vss vss 0.72fF
C19 csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C20 csvco_branch_2/cap_vco_0/t vss 7.10fF
C21 csvco_branch_2/inverter_csvco_0/vss vss 0.62fF
C22 csvco_branch_1/in vss 1.58fF
C23 csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C24 out_vco vss 0.67fF
C25 D0 vss -1.55fF
C26 vdd vss 31.40fF
C27 csvco_branch_0/cap_vco_0/t vss 7.10fF
C28 csvco_branch_0/inverter_csvco_0/vss vss 0.66fF
C29 vctrl vss 11.02fF
C30 csvco_branch_2/vbp vss 0.77fF
.ends

.subckt ring_osc_buffer vss in_vco vdd o1 out_div out_pad
Xinverter_min_x4_0 o1 vss out_div vdd inverter_min_x4
Xinverter_min_x4_1 out_div vss out_pad vdd inverter_min_x4
Xinverter_min_x2_0 in_vco o1 vss vdd inverter_min_x2
C0 vdd o1 0.09fF
C1 out_div vdd 0.17fF
C2 out_div out_pad 0.15fF
C3 out_div o1 0.11fF
C4 vdd out_pad 0.10fF
C5 in_vco vss 0.83fF
C6 out_pad vss 0.70fF
C7 out_div vss 3.00fF
C8 vdd vss 14.54fF
C9 o1 vss 2.72fF
.ends

.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X a_194_125# a_355_368# a_455_87#
+ a_158_392#
X0 X B a_455_87# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 X a_194_125# a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_194_125# B a_158_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_158_392# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_355_368# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_194_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 a_455_87# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND B a_194_125# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X9 VGND a_194_125# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
C0 VPB VPWR 0.06fF
C1 B VGND 0.10fF
C2 a_355_368# VPWR 0.37fF
C3 a_355_368# A 0.02fF
C4 B VPWR 0.09fF
C5 a_194_125# X 0.29fF
C6 VGND VPWR 0.01fF
C7 B A 0.28fF
C8 A VGND 0.31fF
C9 A VPWR 0.15fF
C10 a_355_368# a_194_125# 0.51fF
C11 B a_194_125# 0.57fF
C12 a_355_368# X 0.17fF
C13 a_194_125# VGND 0.25fF
C14 a_194_125# a_158_392# 0.06fF
C15 B X 0.13fF
C16 VGND X 0.28fF
C17 a_194_125# VPWR 0.33fF
C18 a_194_125# A 0.18fF
C19 VPWR X 0.07fF
C20 B a_355_368# 0.08fF
C21 VGND VNB 0.78fF
C22 X VNB 0.21fF
C23 VPWR VNB 0.78fF
C24 B VNB 0.56fF
C25 A VNB 0.70fF
C26 VPB VNB 0.77fF
C27 a_355_368# VNB 0.08fF
C28 a_194_125# VNB 0.40fF
.ends

.subckt sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X a_143_136# a_56_136#
X0 VGND B a_143_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 X a_56_136# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VPWR B a_56_136# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_143_136# A a_56_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_56_136# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 X a_56_136# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
C0 A B 0.08fF
C1 A a_56_136# 0.17fF
C2 VPWR B 0.02fF
C3 VPWR a_56_136# 0.57fF
C4 B X 0.02fF
C5 X a_56_136# 0.26fF
C6 A VGND 0.21fF
C7 B a_56_136# 0.30fF
C8 X VGND 0.15fF
C9 VPWR A 0.07fF
C10 VPWR VPB 0.04fF
C11 VPWR X 0.20fF
C12 B VGND 0.03fF
C13 VGND a_56_136# 0.06fF
C14 VGND VNB 0.50fF
C15 X VNB 0.23fF
C16 VPWR VNB 0.50fF
C17 B VNB 0.24fF
C18 A VNB 0.36fF
C19 VPB VNB 0.48fF
C20 a_56_136# VNB 0.38fF
.ends

.subckt sky130_fd_sc_hs__or2_1 A B VGND VNB VPB VPWR X a_152_368# a_63_368#
X0 VPWR A a_152_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_152_368# B a_63_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 X a_63_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 X a_63_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_63_368# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X5 VGND A a_63_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
C0 X VGND 0.16fF
C1 A a_63_368# 0.28fF
C2 VGND B 0.11fF
C3 a_152_368# a_63_368# 0.03fF
C4 a_63_368# VGND 0.27fF
C5 X VPWR 0.18fF
C6 VPWR VPB 0.04fF
C7 VPWR B 0.01fF
C8 X A 0.02fF
C9 VPWR A 0.05fF
C10 A B 0.10fF
C11 X a_63_368# 0.33fF
C12 VPWR a_63_368# 0.29fF
C13 a_63_368# B 0.14fF
C14 VGND VNB 0.53fF
C15 X VNB 0.24fF
C16 A VNB 0.21fF
C17 B VNB 0.31fF
C18 VPWR VNB 0.46fF
C19 VPB VNB 0.48fF
C20 a_63_368# VNB 0.37fF
.ends

.subckt div_by_5 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_1/latch_diff_0/D
+ nCLK DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/D DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in
+ vdd DFlipFlop_2/latch_diff_0/nD Q0 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ CLK DFlipFlop_2/latch_diff_1/D vss DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ sky130_fd_sc_hs__and2_1_0/a_56_136# nQ0 DFlipFlop_1/latch_diff_1/nD CLK_5 DFlipFlop_3/latch_diff_0/nD
+ nQ2 DFlipFlop_0/latch_diff_0/D DFlipFlop_2/latch_diff_1/nD DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_1/latch_diff_1/D Q1 DFlipFlop_2/D DFlipFlop_3/latch_diff_0/D DFlipFlop_1/D
+ sky130_fd_sc_hs__xor2_1_0/a_355_368# DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_3/latch_diff_1/nD DFlipFlop_0/latch_diff_1/D Q1_shift DFlipFlop_0/latch_diff_0/nD
+ DFlipFlop_2/nQ DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop_2/latch_diff_0/D
+ sky130_fd_sc_hs__xor2_1_0/a_158_392# DFlipFlop_3/latch_diff_1/D sky130_fd_sc_hs__or2_1_0/a_63_368#
+ DFlipFlop_1/latch_diff_0/nD sky130_fd_sc_hs__and2_1_1/a_143_136# DFlipFlop_0/Q sky130_fd_sc_hs__and2_1_1/a_56_136#
+ sky130_fd_sc_hs__xor2_1_0/a_194_125# DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ sky130_fd_sc_hs__and2_1_0/a_143_136#
Xsky130_fd_sc_hs__xor2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_2/D sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ sky130_fd_sc_hs__xor2_1_0/a_355_368# sky130_fd_sc_hs__xor2_1_0/a_455_87# sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ sky130_fd_sc_hs__xor2_1
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vss DFlipFlop_0/latch_diff_1/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ nQ2 DFlipFlop_0/Q DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/D DFlipFlop_0/latch_diff_1/m1_657_280#
+ DFlipFlop_0/latch_diff_0/D vdd CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ nCLK DFlipFlop_0/latch_diff_0/nD DFlipFlop
XDFlipFlop_1 DFlipFlop_1/latch_diff_0/m1_657_280# vss DFlipFlop_1/latch_diff_1/D DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in
+ nQ0 Q0 DFlipFlop_1/latch_diff_1/nD DFlipFlop_1/D DFlipFlop_1/latch_diff_1/m1_657_280#
+ DFlipFlop_1/latch_diff_0/D vdd CLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ nCLK DFlipFlop_1/latch_diff_0/nD DFlipFlop
XDFlipFlop_2 DFlipFlop_2/latch_diff_0/m1_657_280# vss DFlipFlop_2/latch_diff_1/D DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_2/nQ Q1 DFlipFlop_2/latch_diff_1/nD DFlipFlop_2/D DFlipFlop_2/latch_diff_1/m1_657_280#
+ DFlipFlop_2/latch_diff_0/D vdd CLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ nCLK DFlipFlop_2/latch_diff_0/nD DFlipFlop
XDFlipFlop_3 DFlipFlop_3/latch_diff_0/m1_657_280# vss DFlipFlop_3/latch_diff_1/D DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_3/nQ Q1_shift DFlipFlop_3/latch_diff_1/nD Q1 DFlipFlop_3/latch_diff_1/m1_657_280#
+ DFlipFlop_3/latch_diff_0/D vdd nCLK DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out
+ CLK DFlipFlop_3/latch_diff_0/nD DFlipFlop
Xsky130_fd_sc_hs__and2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_0/D sky130_fd_sc_hs__and2_1_0/a_143_136#
+ sky130_fd_sc_hs__and2_1_0/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__and2_1_1 nQ2 nQ0 vss vss vdd vdd DFlipFlop_1/D sky130_fd_sc_hs__and2_1_1/a_143_136#
+ sky130_fd_sc_hs__and2_1_1/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__or2_1_0 Q1 Q1_shift vss vss vdd vdd CLK_5 sky130_fd_sc_hs__or2_1_0/a_152_368#
+ sky130_fd_sc_hs__or2_1_0/a_63_368# sky130_fd_sc_hs__or2_1
C0 CLK DFlipFlop_2/latch_diff_1/D 0.14fF
C1 Q1 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in 0.21fF
C2 Q1_shift DFlipFlop_3/nQ 0.04fF
C3 vdd sky130_fd_sc_hs__xor2_1_0/a_355_368# 0.03fF
C4 vdd DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C5 DFlipFlop_1/latch_diff_1/m1_657_280# nQ0 0.21fF
C6 DFlipFlop_0/latch_diff_0/D Q0 0.42fF
C7 sky130_fd_sc_hs__or2_1_0/a_63_368# vdd 0.02fF
C8 nQ0 DFlipFlop_1/latch_diff_1/D 0.91fF
C9 nCLK sky130_fd_sc_hs__xor2_1_0/a_194_125# 0.11fF
C10 DFlipFlop_3/nQ Q1 0.10fF
C11 DFlipFlop_0/D sky130_fd_sc_hs__and2_1_0/a_56_136# 0.04fF
C12 vdd DFlipFlop_2/nQ 0.02fF
C13 CLK DFlipFlop_1/latch_diff_1/D 0.14fF
C14 DFlipFlop_2/D sky130_fd_sc_hs__xor2_1_0/a_194_125# 0.08fF
C15 nCLK Q1 -0.01fF
C16 nCLK nQ2 0.10fF
C17 DFlipFlop_3/latch_diff_1/nD CLK 0.16fF
C18 DFlipFlop_2/D Q1 0.10fF
C19 Q1 sky130_fd_sc_hs__and2_1_0/a_56_136# 0.14fF
C20 DFlipFlop_0/D Q0 0.39fF
C21 CLK DFlipFlop_3/latch_diff_0/D 0.11fF
C22 DFlipFlop_1/latch_diff_1/nD nQ0 0.88fF
C23 nQ0 sky130_fd_sc_hs__and2_1_1/a_56_136# 0.01fF
C24 nCLK DFlipFlop_2/latch_diff_1/m1_657_280# 0.28fF
C25 sky130_fd_sc_hs__xor2_1_0/a_194_125# Q0 0.26fF
C26 DFlipFlop_1/latch_diff_1/nD CLK 0.09fF
C27 CLK sky130_fd_sc_hs__and2_1_1/a_56_136# 0.06fF
C28 vdd DFlipFlop_0/D 0.19fF
C29 Q1_shift vdd 0.10fF
C30 vdd sky130_fd_sc_hs__xor2_1_0/a_194_125# 0.03fF
C31 sky130_fd_sc_hs__or2_1_0/a_63_368# CLK_5 0.06fF
C32 Q1 Q0 9.65fF
C33 Q0 nQ2 0.23fF
C34 vdd Q1 9.49fF
C35 vdd nQ2 0.04fF
C36 Q1 DFlipFlop_2/latch_diff_0/D 0.42fF
C37 CLK DFlipFlop_2/latch_diff_1/nD 0.09fF
C38 DFlipFlop_0/latch_diff_1/nD CLK 0.02fF
C39 nCLK DFlipFlop_3/latch_diff_0/m1_657_280# 0.27fF
C40 CLK nQ0 0.19fF
C41 sky130_fd_sc_hs__and2_1_1/a_143_136# nQ0 0.04fF
C42 DFlipFlop_1/latch_diff_0/D nQ0 0.09fF
C43 DFlipFlop_0/latch_diff_1/D Q0 0.23fF
C44 CLK sky130_fd_sc_hs__and2_1_1/a_143_136# 0.03fF
C45 Q1 DFlipFlop_2/latch_diff_1/D 0.23fF
C46 DFlipFlop_1/D DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C47 nCLK DFlipFlop_0/Q 0.11fF
C48 nCLK DFlipFlop_3/latch_diff_1/D 0.14fF
C49 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_0/D 0.02fF
C50 nCLK DFlipFlop_1/D 0.14fF
C51 Q1 DFlipFlop_3/latch_diff_0/nD 0.08fF
C52 DFlipFlop_1/latch_diff_1/D Q1 -0.10fF
C53 CLK DFlipFlop_2/latch_diff_0/m1_657_280# 0.28fF
C54 sky130_fd_sc_hs__and2_1_0/a_143_136# Q1 0.02fF
C55 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in Q1 0.09fF
C56 nCLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in 0.14fF
C57 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in Q1 0.20fF
C58 DFlipFlop_3/latch_diff_1/nD Q1 1.24fF
C59 DFlipFlop_0/Q Q0 0.21fF
C60 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out CLK -0.31fF
C61 CLK DFlipFlop_2/nQ 0.13fF
C62 DFlipFlop_3/latch_diff_0/D Q1 0.09fF
C63 DFlipFlop_1/D Q0 0.07fF
C64 CLK DFlipFlop_3/latch_diff_1/m1_657_280# 0.27fF
C65 DFlipFlop_1/latch_diff_1/nD Q1 0.10fF
C66 nCLK DFlipFlop_3/nQ 0.02fF
C67 sky130_fd_sc_hs__and2_1_1/a_56_136# nQ2 0.01fF
C68 vdd DFlipFlop_1/D 0.25fF
C69 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in Q0 0.42fF
C70 DFlipFlop_2/D nCLK 0.41fF
C71 Q1_shift sky130_fd_sc_hs__or2_1_0/a_152_368# -0.04fF
C72 Q1 DFlipFlop_2/latch_diff_1/nD 0.21fF
C73 DFlipFlop_0/latch_diff_1/nD Q1 0.10fF
C74 nQ0 Q1 0.06fF
C75 nQ0 nQ2 0.03fF
C76 vdd DFlipFlop_3/nQ 0.02fF
C77 CLK Q1 -0.10fF
C78 nCLK Q0 0.20fF
C79 CLK nQ2 0.17fF
C80 vdd DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out 0.02fF
C81 DFlipFlop_2/D Q0 0.25fF
C82 DFlipFlop_1/latch_diff_0/D Q1 0.18fF
C83 sky130_fd_sc_hs__and2_1_1/a_143_136# nQ2 0.01fF
C84 Q0 sky130_fd_sc_hs__and2_1_0/a_56_136# 0.17fF
C85 vdd nCLK 0.34fF
C86 nCLK DFlipFlop_2/latch_diff_0/D 0.11fF
C87 vdd DFlipFlop_2/D 0.07fF
C88 vdd sky130_fd_sc_hs__and2_1_0/a_56_136# 0.02fF
C89 sky130_fd_sc_hs__or2_1_0/a_63_368# Q1_shift -0.27fF
C90 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out Q1 0.15fF
C91 DFlipFlop_0/latch_diff_1/D CLK 0.03fF
C92 DFlipFlop_0/latch_diff_1/m1_657_280# nQ2 0.05fF
C93 nCLK DFlipFlop_2/latch_diff_1/D 0.08fF
C94 sky130_fd_sc_hs__and2_1_1/a_56_136# DFlipFlop_1/D 0.04fF
C95 sky130_fd_sc_hs__or2_1_0/a_63_368# Q1 0.10fF
C96 vdd DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in 0.03fF
C97 vdd Q0 5.33fF
C98 Q1 DFlipFlop_2/nQ 0.31fF
C99 DFlipFlop_0/latch_diff_0/m1_657_280# CLK 0.28fF
C100 Q1 DFlipFlop_0/latch_diff_0/D 0.15fF
C101 Q1 DFlipFlop_3/latch_diff_1/m1_657_280# 0.28fF
C102 nCLK DFlipFlop_1/latch_diff_1/m1_657_280# 0.28fF
C103 nCLK DFlipFlop_3/latch_diff_0/nD 0.08fF
C104 nCLK DFlipFlop_1/latch_diff_1/D 0.08fF
C105 DFlipFlop_2/D DFlipFlop_1/latch_diff_1/m1_657_280# 0.04fF
C106 nCLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in -0.33fF
C107 nQ0 DFlipFlop_1/D 0.12fF
C108 DFlipFlop_3/latch_diff_1/nD nCLK 0.09fF
C109 CLK DFlipFlop_0/Q 0.08fF
C110 DFlipFlop_3/latch_diff_1/D CLK 0.08fF
C111 DFlipFlop_0/D Q1 0.13fF
C112 CLK DFlipFlop_1/D 0.21fF
C113 Q1_shift Q1 0.36fF
C114 DFlipFlop_1/latch_diff_1/m1_657_280# Q0 0.01fF
C115 DFlipFlop_1/latch_diff_0/nD nQ0 0.08fF
C116 nCLK DFlipFlop_1/latch_diff_1/nD 0.16fF
C117 DFlipFlop_1/latch_diff_1/D Q0 0.06fF
C118 CLK DFlipFlop_1/latch_diff_0/nD 0.08fF
C119 sky130_fd_sc_hs__and2_1_0/a_143_136# Q0 0.03fF
C120 vdd CLK_5 0.15fF
C121 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in Q0 0.33fF
C122 Q1 nQ2 0.07fF
C123 DFlipFlop_1/latch_diff_0/m1_657_280# nQ0 0.25fF
C124 vdd DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.02fF
C125 Q1 DFlipFlop_2/latch_diff_1/m1_657_280# 0.03fF
C126 vdd DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in 0.03fF
C127 CLK DFlipFlop_1/latch_diff_0/m1_657_280# 0.28fF
C128 DFlipFlop_3/nQ CLK 0.01fF
C129 DFlipFlop_1/latch_diff_1/nD Q0 0.21fF
C130 nCLK DFlipFlop_2/latch_diff_1/nD 0.16fF
C131 nCLK DFlipFlop_0/latch_diff_1/nD 0.05fF
C132 CLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out 0.15fF
C133 nCLK nQ0 0.09fF
C134 vdd sky130_fd_sc_hs__and2_1_1/a_56_136# 0.04fF
C135 DFlipFlop_0/latch_diff_1/D Q1 0.06fF
C136 DFlipFlop_2/D CLK 0.14fF
C137 nCLK DFlipFlop_1/latch_diff_0/D 0.11fF
C138 nCLK sky130_fd_sc_hs__xor2_1_0/a_455_87# 0.02fF
C139 DFlipFlop_2/latch_diff_0/nD CLK 0.08fF
C140 DFlipFlop_3/latch_diff_0/m1_657_280# Q1 0.28fF
C141 DFlipFlop_0/latch_diff_1/nD Q0 0.21fF
C142 nQ0 Q0 0.33fF
C143 DFlipFlop_2/D sky130_fd_sc_hs__xor2_1_0/a_455_87# 0.08fF
C144 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in CLK 0.03fF
C145 CLK Q0 0.08fF
C146 nCLK DFlipFlop_0/latch_diff_1/m1_657_280# 0.28fF
C147 nCLK DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out 0.05fF
C148 vdd nQ0 0.11fF
C149 DFlipFlop_1/latch_diff_0/D Q0 0.42fF
C150 vdd CLK 0.41fF
C151 DFlipFlop_0/Q Q1 0.13fF
C152 DFlipFlop_3/latch_diff_1/D Q1 0.79fF
C153 nCLK DFlipFlop_2/nQ 0.09fF
C154 DFlipFlop_0/Q nQ2 0.09fF
C155 Q1 DFlipFlop_1/D 0.03fF
C156 sky130_fd_sc_hs__xor2_1_0/a_355_368# Q0 0.03fF
C157 CLK_5 vss -0.18fF
C158 sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.38fF
C159 sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.41fF
C160 sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C161 DFlipFlop_3/nQ vss 0.52fF
C162 Q1_shift vss -0.29fF
C163 DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.64fF
C164 DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C165 DFlipFlop_3/latch_diff_1/D vss -1.73fF
C166 DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C167 DFlipFlop_3/latch_diff_0/D vss 0.96fF
C168 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.94fF
C169 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.85fF
C170 DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C171 DFlipFlop_2/nQ vss 0.50fF
C172 Q1 vss 8.55fF
C173 DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.72fF
C174 DFlipFlop_2/latch_diff_1/nD vss 0.58fF
C175 DFlipFlop_2/latch_diff_1/D vss -1.72fF
C176 DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C177 DFlipFlop_2/latch_diff_0/D vss 0.96fF
C178 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.89fF
C179 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C180 DFlipFlop_2/D vss 5.34fF
C181 DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C182 nQ0 vss 3.42fF
C183 Q0 vss 0.53fF
C184 DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.62fF
C185 DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C186 DFlipFlop_1/latch_diff_1/D vss -1.73fF
C187 DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C188 DFlipFlop_1/latch_diff_0/D vss 0.96fF
C189 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C190 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.78fF
C191 DFlipFlop_1/D vss 3.72fF
C192 DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C193 nQ2 vss 2.05fF
C194 DFlipFlop_0/Q vss -0.94fF
C195 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.61fF
C196 nCLK vss 0.96fF
C197 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C198 DFlipFlop_0/latch_diff_1/D vss -1.73fF
C199 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C200 CLK vss 0.20fF
C201 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C202 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.88fF
C203 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C204 DFlipFlop_0/D vss 4.04fF
C205 DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C206 vdd vss 146.76fF
C207 sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C208 sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.42fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AZESM8 a_n63_n151# a_n33_n125# a_n255_n151# a_33_n151#
+ a_n225_n125# a_63_n125# a_n129_n125# a_n159_n151# w_n455_n335# a_225_n151# a_255_n125#
+ a_129_n151# a_159_n125# a_n317_n125#
X0 a_159_n125# a_129_n151# a_63_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n225_n125# a_n255_n151# a_n317_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_63_n125# a_33_n151# a_n33_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_n129_n125# a_n159_n151# a_n225_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n33_n125# a_n63_n151# a_n129_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_255_n125# a_225_n151# a_159_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n129_n125# a_63_n125# 0.13fF
C1 a_255_n125# a_n129_n125# 0.06fF
C2 a_n255_n151# a_n159_n151# 0.02fF
C3 a_n33_n125# a_63_n125# 0.36fF
C4 a_255_n125# a_n33_n125# 0.08fF
C5 a_n63_n151# a_n159_n151# 0.02fF
C6 a_n225_n125# a_n317_n125# 0.36fF
C7 a_159_n125# a_n225_n125# 0.06fF
C8 a_255_n125# a_63_n125# 0.13fF
C9 a_n129_n125# a_n225_n125# 0.36fF
C10 a_n129_n125# a_n317_n125# 0.13fF
C11 a_n129_n125# a_159_n125# 0.08fF
C12 a_225_n151# a_129_n151# 0.02fF
C13 a_n33_n125# a_n225_n125# 0.13fF
C14 a_n33_n125# a_n317_n125# 0.08fF
C15 a_n33_n125# a_159_n125# 0.13fF
C16 a_n225_n125# a_63_n125# 0.08fF
C17 a_n129_n125# a_n33_n125# 0.36fF
C18 a_n63_n151# a_33_n151# 0.02fF
C19 a_33_n151# a_129_n151# 0.02fF
C20 a_63_n125# a_n317_n125# 0.06fF
C21 a_159_n125# a_63_n125# 0.36fF
C22 a_255_n125# a_159_n125# 0.36fF
C23 a_255_n125# w_n455_n335# 0.14fF
C24 a_159_n125# w_n455_n335# 0.08fF
C25 a_63_n125# w_n455_n335# 0.07fF
C26 a_n33_n125# w_n455_n335# 0.08fF
C27 a_n129_n125# w_n455_n335# 0.07fF
C28 a_n225_n125# w_n455_n335# 0.08fF
C29 a_n317_n125# w_n455_n335# 0.14fF
C30 a_225_n151# w_n455_n335# 0.05fF
C31 a_129_n151# w_n455_n335# 0.05fF
C32 a_33_n151# w_n455_n335# 0.05fF
C33 a_n63_n151# w_n455_n335# 0.05fF
C34 a_n159_n151# w_n455_n335# 0.05fF
C35 a_n255_n151# w_n455_n335# 0.05fF
.ends

.subckt sky130_fd_pr__pfet_01v8_XJXT7S VSUBS a_n33_n125# a_n255_n154# a_33_n154# a_n225_n125#
+ a_n159_n154# a_63_n125# a_n129_n125# a_225_n154# a_129_n154# a_255_n125# a_159_n125#
+ a_n317_n125# w_n455_n344# a_n63_n154#
X0 a_n129_n125# a_n159_n154# a_n225_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n33_n125# a_n63_n154# a_n129_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_255_n125# a_225_n154# a_159_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_159_n125# a_129_n154# a_63_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n225_n125# a_n255_n154# a_n317_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_63_n125# a_33_n154# a_n33_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 w_n455_n344# a_255_n125# 0.11fF
C1 w_n455_n344# a_159_n125# 0.06fF
C2 a_n225_n125# a_n33_n125# 0.13fF
C3 a_n129_n125# a_63_n125# 0.13fF
C4 a_n255_n154# a_n159_n154# 0.02fF
C5 a_255_n125# a_n33_n125# 0.08fF
C6 a_n129_n125# a_n317_n125# 0.13fF
C7 a_n33_n125# a_159_n125# 0.13fF
C8 a_n129_n125# w_n455_n344# 0.04fF
C9 a_n225_n125# a_159_n125# 0.06fF
C10 a_n129_n125# a_n33_n125# 0.36fF
C11 a_255_n125# a_159_n125# 0.36fF
C12 a_63_n125# a_n317_n125# 0.06fF
C13 a_n129_n125# a_n225_n125# 0.36fF
C14 w_n455_n344# a_63_n125# 0.04fF
C15 a_33_n154# a_129_n154# 0.02fF
C16 w_n455_n344# a_n317_n125# 0.11fF
C17 a_n129_n125# a_255_n125# 0.06fF
C18 a_n129_n125# a_159_n125# 0.08fF
C19 a_63_n125# a_n33_n125# 0.36fF
C20 a_n317_n125# a_n33_n125# 0.08fF
C21 w_n455_n344# a_n33_n125# 0.05fF
C22 a_225_n154# a_129_n154# 0.02fF
C23 a_63_n125# a_n225_n125# 0.08fF
C24 a_n63_n154# a_n159_n154# 0.02fF
C25 a_n317_n125# a_n225_n125# 0.36fF
C26 a_33_n154# a_n63_n154# 0.02fF
C27 w_n455_n344# a_n225_n125# 0.06fF
C28 a_63_n125# a_255_n125# 0.13fF
C29 a_63_n125# a_159_n125# 0.36fF
C30 a_255_n125# VSUBS 0.03fF
C31 a_159_n125# VSUBS 0.03fF
C32 a_63_n125# VSUBS 0.03fF
C33 a_n33_n125# VSUBS 0.03fF
C34 a_n129_n125# VSUBS 0.03fF
C35 a_n225_n125# VSUBS 0.03fF
C36 a_n317_n125# VSUBS 0.03fF
C37 a_225_n154# VSUBS 0.05fF
C38 a_129_n154# VSUBS 0.05fF
C39 a_33_n154# VSUBS 0.05fF
C40 a_n63_n154# VSUBS 0.05fF
C41 a_n159_n154# VSUBS 0.05fF
C42 a_n255_n154# VSUBS 0.05fF
C43 w_n455_n344# VSUBS 2.96fF
.ends

.subckt inverter_cp_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_AZESM8_0 in vss in in vss out out in vss in out in vss out
+ sky130_fd_pr__nfet_01v8_AZESM8
Xsky130_fd_pr__pfet_01v8_XJXT7S_0 vss vdd in in vdd in out out in in out vdd out vdd
+ in sky130_fd_pr__pfet_01v8_XJXT7S
C0 vdd in 0.04fF
C1 in out 0.85fF
C2 vdd out 0.29fF
C3 vdd vss 5.90fF
C4 out vss 1.30fF
C5 in vss 1.82fF
.ends

.subckt pfd_cp_interface vss inverter_cp_x1_2/in vdd inverter_cp_x1_0/out Down QA
+ QB nDown Up nUp
Xinverter_cp_x2_0 nDown Down vss vdd inverter_cp_x2
Xinverter_cp_x2_1 Up nUp vss vdd inverter_cp_x2
Xtrans_gate_0 nDown inverter_cp_x1_0/out vss vdd trans_gate
Xinverter_cp_x1_0 inverter_cp_x1_0/out QB vss vdd inverter_cp_x1
Xinverter_cp_x1_2 Up inverter_cp_x1_2/in vss vdd inverter_cp_x1
Xinverter_cp_x1_1 inverter_cp_x1_2/in QA vss vdd inverter_cp_x1
C0 Up inverter_cp_x1_2/in 0.12fF
C1 Down vdd 0.09fF
C2 nUp vdd 0.14fF
C3 Down inverter_cp_x1_0/out 0.12fF
C4 vdd QA 0.02fF
C5 Down nDown 0.23fF
C6 vdd inverter_cp_x1_0/out 0.25fF
C7 nDown vdd 0.80fF
C8 QB vdd 0.02fF
C9 nDown inverter_cp_x1_0/out 0.11fF
C10 nUp Up 0.20fF
C11 Up vdd 0.60fF
C12 vdd inverter_cp_x1_2/in 0.42fF
C13 inverter_cp_x1_2/in vss 2.01fF
C14 QA vss 1.09fF
C15 inverter_cp_x1_0/out vss 2.00fF
C16 QB vss 1.09fF
C17 vdd vss 28.96fF
C18 nUp vss 1.32fF
C19 Up vss 2.53fF
C20 Down vss 1.26fF
C21 nDown vss 2.98fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4F35BC VSUBS a_n129_n90# w_n359_n309# a_n63_n116#
+ a_n159_n207# a_63_n90# a_n33_n90# a_n221_n90# a_159_n90#
X0 a_159_n90# a_n63_n116# a_63_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n129_n90# a_n159_n207# a_n221_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X2 a_63_n90# a_n159_n207# a_n33_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3 a_n33_n90# a_n63_n116# a_n129_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_n63_n116# a_n159_n207# 0.12fF
C1 w_n359_n309# a_63_n90# 0.06fF
C2 w_n359_n309# a_n221_n90# 0.09fF
C3 a_63_n90# a_n129_n90# 0.09fF
C4 a_n33_n90# w_n359_n309# 0.05fF
C5 w_n359_n309# a_159_n90# 0.09fF
C6 a_n221_n90# a_n129_n90# 0.26fF
C7 a_n33_n90# a_n129_n90# 0.26fF
C8 a_n129_n90# a_159_n90# 0.06fF
C9 a_63_n90# a_n221_n90# 0.06fF
C10 a_n33_n90# a_63_n90# 0.26fF
C11 a_63_n90# a_159_n90# 0.26fF
C12 a_n33_n90# a_n221_n90# 0.09fF
C13 a_n221_n90# a_159_n90# 0.04fF
C14 a_n33_n90# a_159_n90# 0.09fF
C15 w_n359_n309# a_n129_n90# 0.06fF
C16 a_159_n90# VSUBS 0.03fF
C17 a_63_n90# VSUBS 0.03fF
C18 a_n33_n90# VSUBS 0.03fF
C19 a_n129_n90# VSUBS 0.03fF
C20 a_n221_n90# VSUBS 0.03fF
C21 a_n159_n207# VSUBS 0.30fF
C22 a_n63_n116# VSUBS 0.37fF
C23 w_n359_n309# VSUBS 2.23fF
.ends

.subckt sky130_fd_pr__nfet_01v8_C3YG4M a_n33_n45# a_33_n71# a_n129_71# w_n263_n255#
+ a_n125_n45# a_63_n45#
X0 a_63_n45# a_33_n71# a_n33_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n129_71# a_n125_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_63_n45# a_n33_n45# 0.13fF
C1 a_n129_71# a_33_n71# 0.04fF
C2 a_63_n45# a_n125_n45# 0.05fF
C3 a_n33_n45# a_n125_n45# 0.13fF
C4 a_63_n45# w_n263_n255# 0.04fF
C5 a_n33_n45# w_n263_n255# 0.04fF
C6 a_n125_n45# w_n263_n255# 0.04fF
C7 a_33_n71# w_n263_n255# 0.11fF
C8 a_n129_71# w_n263_n255# 0.14fF
.ends

.subckt nor_pfd sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd A B
Xsky130_fd_pr__pfet_01v8_4F35BC_0 vss sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vdd B A sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out vdd vdd sky130_fd_pr__pfet_01v8_4F35BC
Xsky130_fd_pr__nfet_01v8_C3YG4M_0 out B A vss vss vss sky130_fd_pr__nfet_01v8_C3YG4M
C0 vdd sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.02fF
C1 out sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.08fF
C2 out vdd 0.11fF
C3 vdd A 0.09fF
C4 out A 0.06fF
C5 sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vdd 0.02fF
C6 out B 0.40fF
C7 A B 0.24fF
C8 sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C9 out vss 0.45fF
C10 sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C11 A vss 0.83fF
C12 B vss 1.09fF
C13 vdd vss 3.79fF
.ends

.subckt dff_pfd vss vdd nor_pfd_2/A Q CLK nor_pfd_3/A nor_pfd_2/B Reset
Xnor_pfd_0 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_2/A nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd CLK Q nor_pfd
Xnor_pfd_1 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# Q nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd nor_pfd_2/A nor_pfd_3/A nor_pfd
Xnor_pfd_2 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_3/A nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd nor_pfd_2/A nor_pfd_2/B nor_pfd
Xnor_pfd_3 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_2/B nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd nor_pfd_3/A Reset nor_pfd
C0 Reset nor_pfd_3/A 0.12fF
C1 vdd nor_pfd_2/A -0.01fF
C2 CLK Q 0.04fF
C3 Reset Q 0.14fF
C4 nor_pfd_3/A Q 0.98fF
C5 vdd nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.06fF
C6 vdd nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.06fF
C7 nor_pfd_3/A nor_pfd_2/A 0.38fF
C8 vdd nor_pfd_2/B 0.02fF
C9 nor_pfd_2/A Q 1.38fF
C10 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vdd 0.06fF
C11 nor_pfd_2/B Reset 0.43fF
C12 nor_pfd_2/B nor_pfd_3/A 0.58fF
C13 vdd nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.06fF
C14 nor_pfd_2/B Q 2.22fF
C15 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vdd 0.06fF
C16 vdd nor_pfd_3/A 0.09fF
C17 vdd nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.06fF
C18 vdd Q 0.08fF
C19 nor_pfd_2/B nor_pfd_2/A 0.05fF
C20 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C21 nor_pfd_2/B vss 1.42fF
C22 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C23 nor_pfd_3/A vss 3.16fF
C24 Reset vss 1.48fF
C25 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C26 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C27 nor_pfd_2/A vss 2.56fF
C28 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C29 Q vss 2.77fF
C30 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C31 vdd vss 16.42fF
C32 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C33 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C34 CLK vss 0.95fF
.ends

.subckt sky130_fd_pr__nfet_01v8_ZCYAJJ w_n359_n255# a_n33_n45# a_n159_n173# a_n221_n45#
+ a_159_n45# a_n63_n71# a_n129_n45# a_63_n45#
X0 a_63_n45# a_n159_n173# a_n33_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n63_n71# a_n129_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X2 a_159_n45# a_n63_n71# a_63_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X3 a_n129_n45# a_n159_n173# a_n221_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_159_n45# a_n221_n45# 0.02fF
C1 a_63_n45# a_n221_n45# 0.03fF
C2 a_n221_n45# a_n129_n45# 0.13fF
C3 a_n63_n71# a_n159_n173# 0.10fF
C4 a_63_n45# a_159_n45# 0.13fF
C5 a_159_n45# a_n129_n45# 0.03fF
C6 a_63_n45# a_n129_n45# 0.05fF
C7 a_n33_n45# a_n221_n45# 0.05fF
C8 a_159_n45# a_n33_n45# 0.05fF
C9 a_63_n45# a_n33_n45# 0.13fF
C10 a_n33_n45# a_n129_n45# 0.13fF
C11 a_159_n45# w_n359_n255# 0.04fF
C12 a_63_n45# w_n359_n255# 0.05fF
C13 a_n33_n45# w_n359_n255# 0.05fF
C14 a_n129_n45# w_n359_n255# 0.05fF
C15 a_n221_n45# w_n359_n255# 0.08fF
C16 a_n159_n173# w_n359_n255# 0.31fF
C17 a_n63_n71# w_n359_n255# 0.31fF
.ends

.subckt sky130_fd_pr__pfet_01v8_7T83YG VSUBS a_n125_n90# a_63_n90# a_33_n187# a_n99_n187#
+ a_n33_n90# w_n263_n309#
X0 a_63_n90# a_33_n187# a_n33_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n33_n90# a_n99_n187# a_n125_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_n33_n90# a_n125_n90# 0.26fF
C1 a_63_n90# a_n125_n90# 0.09fF
C2 a_n99_n187# a_33_n187# 0.04fF
C3 a_63_n90# a_n33_n90# 0.26fF
C4 a_63_n90# VSUBS 0.03fF
C5 a_n33_n90# VSUBS 0.03fF
C6 a_n125_n90# VSUBS 0.03fF
C7 a_33_n187# VSUBS 0.12fF
C8 a_n99_n187# VSUBS 0.12fF
C9 w_n263_n309# VSUBS 1.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_ZXAV3F a_n73_n45# a_n33_67# a_15_n45# w_n211_n255#
X0 a_15_n45# a_n33_67# a_n73_n45# w_n211_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_n73_n45# a_15_n45# 0.16fF
C1 a_15_n45# w_n211_n255# 0.08fF
C2 a_n73_n45# w_n211_n255# 0.06fF
C3 a_n33_67# w_n211_n255# 0.10fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4F7GBC VSUBS a_n51_n187# a_n73_n90# a_15_n90# w_n211_n309#
X0 a_15_n90# a_n51_n187# a_n73_n90# w_n211_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_n73_n90# a_15_n90# 0.31fF
C1 a_n73_n90# w_n211_n309# 0.04fF
C2 a_15_n90# w_n211_n309# 0.09fF
C3 a_15_n90# VSUBS 0.03fF
C4 a_n73_n90# VSUBS 0.03fF
C5 a_n51_n187# VSUBS 0.12fF
C6 w_n211_n309# VSUBS 1.24fF
.ends

.subckt and_pfd a_656_410# vss out vdd A B
Xsky130_fd_pr__nfet_01v8_ZCYAJJ_0 vss a_656_410# A vss vss B sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45#
+ sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# sky130_fd_pr__nfet_01v8_ZCYAJJ
Xsky130_fd_pr__pfet_01v8_7T83YG_0 vss vdd vdd B A a_656_410# vdd sky130_fd_pr__pfet_01v8_7T83YG
Xsky130_fd_pr__nfet_01v8_ZXAV3F_0 vss a_656_410# out vss sky130_fd_pr__nfet_01v8_ZXAV3F
Xsky130_fd_pr__pfet_01v8_4F7GBC_0 vss a_656_410# vdd out vdd sky130_fd_pr__pfet_01v8_4F7GBC
C0 a_656_410# out 0.20fF
C1 A vdd 0.05fF
C2 a_656_410# vdd 0.20fF
C3 A B 0.33fF
C4 a_656_410# B 0.30fF
C5 a_656_410# sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# 0.07fF
C6 vdd out 0.10fF
C7 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# B 0.02fF
C8 A a_656_410# 0.04fF
C9 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# out 0.03fF
C10 vdd vss 4.85fF
C11 out vss 0.47fF
C12 a_656_410# vss 1.00fF
C13 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.13fF
C14 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.10fF
C15 A vss 0.85fF
C16 B vss 0.95fF
.ends

.subckt PFD vss vdd Down Up A B Reset
Xdff_pfd_0 vss vdd dff_pfd_0/nor_pfd_2/A Up A dff_pfd_0/nor_pfd_3/A dff_pfd_0/nor_pfd_2/B
+ Reset dff_pfd
Xdff_pfd_1 vss vdd dff_pfd_1/nor_pfd_2/A Down B dff_pfd_1/nor_pfd_3/A dff_pfd_1/nor_pfd_2/B
+ Reset dff_pfd
Xand_pfd_0 and_pfd_0/a_656_410# vss Reset vdd Up Down and_pfd
C0 dff_pfd_1/nor_pfd_2/B vdd 0.04fF
C1 Reset vdd 0.02fF
C2 dff_pfd_0/nor_pfd_2/A vdd 0.13fF
C3 Up Down 0.06fF
C4 dff_pfd_0/nor_pfd_3/A vdd 0.08fF
C5 vdd Down 0.08fF
C6 vdd Up 1.62fF
C7 dff_pfd_1/nor_pfd_3/A vdd 0.08fF
C8 vdd dff_pfd_1/nor_pfd_2/A 0.13fF
C9 vdd dff_pfd_0/nor_pfd_2/B 0.11fF
C10 and_pfd_0/a_656_410# vss 0.99fF
C11 and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C12 and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.05fF
C13 dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C14 dff_pfd_1/nor_pfd_2/B vss 1.51fF
C15 dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C16 dff_pfd_1/nor_pfd_3/A vss 3.14fF
C17 dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C18 dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C19 dff_pfd_1/nor_pfd_2/A vss 2.56fF
C20 dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C21 Down vss 3.74fF
C22 dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C23 vdd vss 44.73fF
C24 dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C25 dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C26 B vss 1.07fF
C27 dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C28 dff_pfd_0/nor_pfd_2/B vss 1.40fF
C29 dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C30 dff_pfd_0/nor_pfd_3/A vss 3.14fF
C31 Reset vss 3.85fF
C32 dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C33 dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C34 dff_pfd_0/nor_pfd_2/A vss 2.56fF
C35 dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C36 Up vss 3.18fF
C37 dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C38 dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C39 dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C40 A vss 1.07fF
.ends


* Top level circuit top_pll_v1

Xloop_filter_0 lf_vc vco_vctrl vss loop_filter
Xcharge_pump_0 nswitch vdd nUp vss Down biasp vco_vctrl pswitch iref_cp nDown Up charge_pump
Xdiv_by_2_0 vss vdd div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in out_by_2 n_out_by_2
+ out_buffer_div_2 out_to_div out_div_2 n_out_buffer_div_2 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out
+ n_out_div_2 div_by_2
Xbuffer_salida_0 buffer_salida_0/a_678_n100# out_to_pad out_to_buffer vss vdd buffer_salida
Xring_osc_0 vco_vctrl vdd vss ring_osc_0/csvco_branch_0/inverter_csvco_0/vss ring_osc_0/csvco_branch_2/vbp
+ vco_D0 ring_osc_0/csvco_branch_2/cap_vco_0/t vco_out ring_osc
Xring_osc_buffer_0 vss vco_out vdd out_first_buffer out_to_div out_to_buffer ring_osc_buffer
Xdiv_by_5_0 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/DFlipFlop_1/latch_diff_0/D
+ n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/nD div_by_5_0/DFlipFlop_0/D div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in
+ vdd div_by_5_0/DFlipFlop_2/latch_diff_0/nD div_5_Q0 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# div_5_nQ0 div_by_5_0/DFlipFlop_1/latch_diff_1/nD
+ out_div_by_5 div_by_5_0/DFlipFlop_3/latch_diff_0/nD div_5_nQ2 div_by_5_0/DFlipFlop_0/latch_diff_0/D
+ div_by_5_0/DFlipFlop_2/latch_diff_1/nD div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_1/latch_diff_1/D div_5_Q1 div_by_5_0/DFlipFlop_2/D div_by_5_0/DFlipFlop_3/latch_diff_0/D
+ div_by_5_0/DFlipFlop_1/D div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_3/latch_diff_1/nD div_by_5_0/DFlipFlop_0/latch_diff_1/D div_5_Q1_shift
+ div_by_5_0/DFlipFlop_0/latch_diff_0/nD div_by_5_0/DFlipFlop_2/nQ div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_2/latch_diff_0/D div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ div_by_5_0/DFlipFlop_3/latch_diff_1/D div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368#
+ div_by_5_0/DFlipFlop_1/latch_diff_0/nD div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136#
+ div_by_5_0/DFlipFlop_0/Q div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136#
+ div_by_5
Xpfd_cp_interface_0 vss pfd_cp_interface_0/inverter_cp_x1_2/in vdd pfd_cp_interface_0/inverter_cp_x1_0/out
+ Down QA QB nDown Up nUp pfd_cp_interface
XPFD_0 vss vdd QB QA in_ref out_div_by_5 pfd_reset PFD
C0 vdd n_out_by_2 1.03fF
C1 div_5_nQ2 n_out_by_2 0.10fF
C2 div_by_5_0/DFlipFlop_2/nQ n_out_by_2 0.10fF
C3 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out out_by_2 0.28fF
C4 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in out_by_2 -0.22fF
C5 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# n_out_by_2 0.12fF
C6 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vdd 0.03fF
C7 div_by_5_0/DFlipFlop_3/latch_diff_1/D out_by_2 0.09fF
C8 n_out_by_2 div_by_5_0/DFlipFlop_0/Q -0.23fF
C9 div_by_5_0/DFlipFlop_1/latch_diff_1/nD out_by_2 0.09fF
C10 div_by_5_0/DFlipFlop_0/D n_out_by_2 -1.48fF
C11 div_by_5_0/DFlipFlop_2/latch_diff_0/nD out_by_2 0.10fF
C12 div_by_5_0/DFlipFlop_1/D n_out_by_2 0.22fF
C13 div_by_5_0/DFlipFlop_0/latch_diff_1/nD out_by_2 0.17fF
C14 vdd Up 0.28fF
C15 nUp vco_vctrl 0.02fF
C16 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# out_div_by_5 0.18fF
C17 vdd iref_cp 0.15fF
C18 nswitch vco_vctrl -0.06fF
C19 biasp nDown 0.26fF
C20 nUp biasp -0.17fF
C21 out_to_buffer out_to_div 0.13fF
C22 nUp nDown -0.09fF
C23 vco_vctrl out_by_2 0.53fF
C24 nswitch nDown 0.76fF
C25 div_by_5_0/DFlipFlop_1/latch_diff_0/nD out_by_2 0.10fF
C26 n_out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/nD 0.10fF
C27 div_5_Q0 n_out_by_2 -0.12fF
C28 Up pswitch 1.98fF
C29 QA vdd -0.04fF
C30 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in n_out_by_2 0.27fF
C31 vco_D0 vdd 0.03fF
C32 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# n_out_by_2 0.02fF
C33 biasp Down 1.24fF
C34 vco_vctrl ring_osc_0/csvco_branch_2/vbp 0.26fF
C35 Down nDown 2.55fF
C36 nswitch Down 0.54fF
C37 div_5_Q1 out_div_by_5 0.01fF
C38 div_by_5_0/DFlipFlop_3/latch_diff_0/D out_by_2 0.11fF
C39 div_5_Q1 vco_vctrl 0.14fF
C40 out_to_div vdd 0.21fF
C41 div_by_5_0/DFlipFlop_3/latch_diff_1/D n_out_by_2 0.24fF
C42 div_by_5_0/DFlipFlop_2/latch_diff_1/D out_by_2 0.23fF
C43 div_by_5_0/DFlipFlop_1/latch_diff_1/nD n_out_by_2 0.24fF
C44 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# out_by_2 0.10fF
C45 div_5_nQ0 out_by_2 0.32fF
C46 div_5_Q1 out_by_2 0.42fF
C47 n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_0/D 0.24fF
C48 div_by_5_0/DFlipFlop_0/latch_diff_1/nD n_out_by_2 0.33fF
C49 out_by_2 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out -0.04fF
C50 div_by_5_0/DFlipFlop_1/latch_diff_1/D out_by_2 0.23fF
C51 vco_vctrl n_out_by_2 0.52fF
C52 div_by_5_0/DFlipFlop_2/latch_diff_1/nD out_by_2 0.09fF
C53 div_by_5_0/DFlipFlop_0/latch_diff_1/D out_by_2 0.33fF
C54 vdd out_div_by_5 0.28fF
C55 vdd vco_vctrl -1.02fF
C56 div_by_5_0/DFlipFlop_0/latch_diff_0/nD out_by_2 0.17fF
C57 div_by_5_0/DFlipFlop_2/D out_by_2 0.22fF
C58 out_to_buffer buffer_salida_0/a_678_n100# 0.22fF
C59 div_5_Q1_shift out_div_by_5 0.05fF
C60 out_to_div div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in -0.16fF
C61 nUp vdd 0.05fF
C62 vdd nDown 0.22fF
C63 div_by_5_0/DFlipFlop_1/latch_diff_0/D n_out_by_2 0.12fF
C64 div_5_nQ2 out_by_2 0.16fF
C65 vdd out_by_2 0.97fF
C66 div_by_5_0/DFlipFlop_2/nQ out_by_2 0.23fF
C67 lf_vc vdd 0.02fF
C68 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392# n_out_by_2 0.01fF
C69 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vco_vctrl -0.36fF
C70 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136# out_by_2 -0.02fF
C71 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out out_by_2 0.09fF
C72 pswitch nDown 0.53fF
C73 nUp pswitch 0.85fF
C74 n_out_by_2 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in -0.20fF
C75 vdd pfd_cp_interface_0/inverter_cp_x1_2/in 0.01fF
C76 out_first_buffer ring_osc_0/csvco_branch_2/cap_vco_0/t 0.03fF
C77 div_by_5_0/DFlipFlop_3/latch_diff_0/nD n_out_by_2 0.11fF
C78 div_by_5_0/DFlipFlop_2/latch_diff_0/D n_out_by_2 0.12fF
C79 n_out_by_2 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in -0.51fF
C80 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out n_out_by_2 -0.11fF
C81 vdd ring_osc_0/csvco_branch_2/vbp 0.03fF
C82 div_by_5_0/DFlipFlop_2/latch_diff_1/D n_out_by_2 0.10fF
C83 vdd ring_osc_0/csvco_branch_2/cap_vco_0/t 0.02fF
C84 div_by_5_0/DFlipFlop_0/D vco_vctrl -0.45fF
C85 vdd div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out 0.04fF
C86 div_5_nQ0 n_out_by_2 0.10fF
C87 biasp Up 0.26fF
C88 div_by_5_0/DFlipFlop_0/Q out_by_2 0.09fF
C89 div_5_Q1 n_out_by_2 1.04fF
C90 vdd buffer_salida_0/a_678_n100# 0.24fF
C91 ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vco_vctrl 0.04fF
C92 nUp Up 2.72fF
C93 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# -0.05fF
C94 out_to_buffer vdd 0.07fF
C95 div_by_5_0/DFlipFlop_0/D out_by_2 0.35fF
C96 div_by_5_0/DFlipFlop_1/D out_by_2 0.38fF
C97 out_to_div div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out -0.12fF
C98 div_5_Q0 vco_vctrl 0.48fF
C99 div_by_5_0/DFlipFlop_1/latch_diff_1/D n_out_by_2 0.10fF
C100 n_out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/nD 0.24fF
C101 div_by_5_0/DFlipFlop_0/latch_diff_1/D n_out_by_2 0.17fF
C102 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# n_out_by_2 0.03fF
C103 div_by_5_0/DFlipFlop_3/latch_diff_1/nD out_by_2 0.23fF
C104 div_5_Q0 out_by_2 0.09fF
C105 iref_cp Down 0.09fF
C106 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# vco_vctrl -0.11fF
C107 div_by_5_0/DFlipFlop_2/D n_out_by_2 0.19fF
C108 PFD_0/and_pfd_0/a_656_410# vss 0.96fF
C109 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C110 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.07fF
C111 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C112 PFD_0/dff_pfd_1/nor_pfd_2/B vss 1.40fF
C113 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C114 PFD_0/dff_pfd_1/nor_pfd_3/A vss 3.14fF
C115 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C116 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C117 PFD_0/dff_pfd_1/nor_pfd_2/A vss 2.55fF
C118 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C119 QB vss 4.46fF
C120 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C121 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C122 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C123 out_div_by_5 vss -0.40fF
C124 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C125 PFD_0/dff_pfd_0/nor_pfd_2/B vss 1.40fF
C126 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C127 PFD_0/dff_pfd_0/nor_pfd_3/A vss 3.14fF
C128 pfd_reset vss 2.17fF
C129 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C130 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C131 PFD_0/dff_pfd_0/nor_pfd_2/A vss 2.55fF
C132 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C133 QA vss 4.31fF
C134 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C135 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C136 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C137 in_ref vss 1.19fF
C138 pfd_cp_interface_0/inverter_cp_x1_2/in vss 1.85fF
C139 pfd_cp_interface_0/inverter_cp_x1_0/out vss 1.87fF
C140 nUp vss 5.50fF
C141 Up vss 2.37fF
C142 Down vss 7.92fF
C143 nDown vss -2.20fF
C144 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C145 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.38fF
C146 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.41fF
C147 div_by_5_0/DFlipFlop_3/nQ vss 0.48fF
C148 div_5_Q1_shift vss -0.14fF
C149 div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.57fF
C150 div_by_5_0/DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C151 div_by_5_0/DFlipFlop_3/latch_diff_1/D vss -1.73fF
C152 div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C153 div_by_5_0/DFlipFlop_3/latch_diff_0/D vss 0.96fF
C154 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C155 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C156 div_by_5_0/DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C157 div_by_5_0/DFlipFlop_2/nQ vss 0.48fF
C158 div_5_Q1 vss 4.28fF
C159 div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C160 div_by_5_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C161 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C162 div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C163 div_by_5_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C164 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C165 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C166 div_by_5_0/DFlipFlop_2/D vss 3.13fF
C167 div_by_5_0/DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C168 div_5_nQ0 vss 0.59fF
C169 div_5_Q0 vss 0.01fF
C170 div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C171 div_by_5_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C172 div_by_5_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C173 div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C174 div_by_5_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C175 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C176 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C177 div_by_5_0/DFlipFlop_1/D vss 3.64fF
C178 div_by_5_0/DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C179 div_5_nQ2 vss 1.24fF
C180 div_by_5_0/DFlipFlop_0/Q vss -0.94fF
C181 div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C182 n_out_by_2 vss -2.62fF
C183 div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C184 div_by_5_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C185 div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C186 out_by_2 vss -4.51fF
C187 div_by_5_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C188 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C189 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C190 div_by_5_0/DFlipFlop_0/D vss 3.96fF
C191 div_by_5_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C192 vdd vss 366.82fF
C193 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C194 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.40fF
C195 out_to_buffer vss 1.57fF
C196 out_to_div vss 4.46fF
C197 out_first_buffer vss 2.88fF
C198 ring_osc_0/csvco_branch_2/in vss 1.60fF
C199 ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C200 ring_osc_0/csvco_branch_1/cap_vco_0/t vss 7.10fF
C201 ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vss 0.52fF
C202 ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C203 ring_osc_0/csvco_branch_2/cap_vco_0/t vss 7.10fF
C204 ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vss 0.52fF
C205 ring_osc_0/csvco_branch_1/in vss 1.58fF
C206 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C207 vco_out vss 1.01fF
C208 vco_D0 vss -4.63fF
C209 ring_osc_0/csvco_branch_0/cap_vco_0/t vss 7.10fF
C210 ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vss 0.52fF
C211 ring_osc_0/csvco_branch_2/vbp vss 0.38fF
C212 out_to_pad vss 7.50fF
C213 buffer_salida_0/a_3996_n100# vss 48.29fF
C214 buffer_salida_0/a_678_n100# vss 13.38fF
C215 n_out_buffer_div_2 vss 1.63fF
C216 out_buffer_div_2 vss 1.60fF
C217 div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C218 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C219 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.89fF
C220 div_by_2_0/DFlipFlop_0/nCLK vss 1.03fF
C221 out_div_2 vss -1.30fF
C222 div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C223 div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C224 div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C225 div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C226 div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C227 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C228 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C229 n_out_div_2 vss 1.95fF
C230 div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C231 nswitch vss 3.73fF
C232 biasp vss 5.44fF
C233 iref_cp vss 2.81fF
C234 vco_vctrl vss -19.28fF
C235 pswitch vss 3.57fF
C236 lf_vc vss -59.89fF
C237 loop_filter_0/res_loop_filter_2/out vss 7.90fF
.end

