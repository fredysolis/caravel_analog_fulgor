**.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
*+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3],wbs_sel_i[2],wbs_sel_i[1],wbs_sel_i[0]
*+ wbs_dat_i[31],wbs_dat_i[30],wbs_dat_i[29],wbs_dat_i[28],wbs_dat_i[27],wbs_dat_i[26],wbs_dat_i[25],wbs_dat_i[24],wbs_dat_i[23],wbs_dat_i[22],wbs_dat_i[21],wbs_dat_i[20],wbs_dat_i[19],wbs_dat_i[18],wbs_dat_i[17],wbs_dat_i[16],wbs_dat_i[15],wbs_dat_i[14],wbs_dat_i[13],wbs_dat_i[12],wbs_dat_i[11],wbs_dat_i[10],wbs_dat_i[9],wbs_dat_i[8],wbs_dat_i[7],wbs_dat_i[6],wbs_dat_i[5],wbs_dat_i[4],wbs_dat_i[3],wbs_dat_i[2],wbs_dat_i[1],wbs_dat_i[0]
*+ wbs_adr_i[31],wbs_adr_i[30],wbs_adr_i[29],wbs_adr_i[28],wbs_adr_i[27],wbs_adr_i[26],wbs_adr_i[25],wbs_adr_i[24],wbs_adr_i[23],wbs_adr_i[22],wbs_adr_i[21],wbs_adr_i[20],wbs_adr_i[19],wbs_adr_i[18],wbs_adr_i[17],wbs_adr_i[16],wbs_adr_i[15],wbs_adr_i[14],wbs_adr_i[13],wbs_adr_i[12],wbs_adr_i[11],wbs_adr_i[10],wbs_adr_i[9],wbs_adr_i[8],wbs_adr_i[7],wbs_adr_i[6],wbs_adr_i[5],wbs_adr_i[4],wbs_adr_i[3],wbs_adr_i[2],wbs_adr_i[1],wbs_adr_i[0] wbs_ack_o
*+ wbs_dat_o[31],wbs_dat_o[30],wbs_dat_o[29],wbs_dat_o[28],wbs_dat_o[27],wbs_dat_o[26],wbs_dat_o[25],wbs_dat_o[24],wbs_dat_o[23],wbs_dat_o[22],wbs_dat_o[21],wbs_dat_o[20],wbs_dat_o[19],wbs_dat_o[18],wbs_dat_o[17],wbs_dat_o[16],wbs_dat_o[15],wbs_dat_o[14],wbs_dat_o[13],wbs_dat_o[12],wbs_dat_o[11],wbs_dat_o[10],wbs_dat_o[9],wbs_dat_o[8],wbs_dat_o[7],wbs_dat_o[6],wbs_dat_o[5],wbs_dat_o[4],wbs_dat_o[3],wbs_dat_o[2],wbs_dat_o[1],wbs_dat_o[0]
*+ la_data_in[127],la_data_in[126],la_data_in[125],la_data_in[124],la_data_in[123],la_data_in[122],la_data_in[121],la_data_in[120],la_data_in[119],la_data_in[118],la_data_in[117],la_data_in[116],la_data_in[115],la_data_in[114],la_data_in[113],la_data_in[112],la_data_in[111],la_data_in[110],la_data_in[109],la_data_in[108],la_data_in[107],la_data_in[106],la_data_in[105],la_data_in[104],la_data_in[103],la_data_in[102],la_data_in[101],la_data_in[100],la_data_in[99],la_data_in[98],la_data_in[97],la_data_in[96],la_data_in[95],la_data_in[94],la_data_in[93],la_data_in[92],la_data_in[91],la_data_in[90],la_data_in[89],la_data_in[88],la_data_in[87],la_data_in[86],la_data_in[85],la_data_in[84],la_data_in[83],la_data_in[82],la_data_in[81],la_data_in[80],la_data_in[79],la_data_in[78],la_data_in[77],la_data_in[76],la_data_in[75],la_data_in[74],la_data_in[73],la_data_in[72],la_data_in[71],la_data_in[70],la_data_in[69],la_data_in[68],la_data_in[67],la_data_in[66],la_data_in[65],la_data_in[64],la_data_in[63],la_data_in[62],la_data_in[61],la_data_in[60],la_data_in[59],la_data_in[58],la_data_in[57],la_data_in[56],la_data_in[55],la_data_in[54],la_data_in[53],la_data_in[52],la_data_in[51],la_data_in[50],la_data_in[49],la_data_in[48],la_data_in[47],la_data_in[46],la_data_in[45],la_data_in[44],la_data_in[43],la_data_in[42],la_data_in[41],la_data_in[40],la_data_in[39],la_data_in[38],la_data_in[37],la_data_in[36],la_data_in[35],la_data_in[34],la_data_in[33],la_data_in[32],la_data_in[31],la_data_in[30],la_data_in[29],la_data_in[28],la_data_in[27],la_data_in[26],la_data_in[25],la_data_in[24],la_data_in[23],la_data_in[22],la_data_in[21],la_data_in[20],la_data_in[19],la_data_in[18],la_data_in[17],la_data_in[16],la_data_in[15],la_data_in[14],la_data_in[13],la_data_in[12],la_data_in[11],la_data_in[10],la_data_in[9],la_data_in[8],la_data_in[7],la_data_in[6],la_data_in[5],la_data_in[4],la_data_in[3],la_data_in[2],la_data_in[1],la_data_in[0]
*+ la_data_out[127],la_data_out[126],la_data_out[125],la_data_out[124],la_data_out[123],la_data_out[122],la_data_out[121],la_data_out[120],la_data_out[119],la_data_out[118],la_data_out[117],la_data_out[116],la_data_out[115],la_data_out[114],la_data_out[113],la_data_out[112],la_data_out[111],la_data_out[110],la_data_out[109],la_data_out[108],la_data_out[107],la_data_out[106],la_data_out[105],la_data_out[104],la_data_out[103],la_data_out[102],la_data_out[101],la_data_out[100],la_data_out[99],la_data_out[98],la_data_out[97],la_data_out[96],la_data_out[95],la_data_out[94],la_data_out[93],la_data_out[92],la_data_out[91],la_data_out[90],la_data_out[89],la_data_out[88],la_data_out[87],la_data_out[86],la_data_out[85],la_data_out[84],la_data_out[83],la_data_out[82],la_data_out[81],la_data_out[80],la_data_out[79],la_data_out[78],la_data_out[77],la_data_out[76],la_data_out[75],la_data_out[74],la_data_out[73],la_data_out[72],la_data_out[71],la_data_out[70],la_data_out[69],la_data_out[68],la_data_out[67],la_data_out[66],la_data_out[65],la_data_out[64],la_data_out[63],la_data_out[62],la_data_out[61],la_data_out[60],la_data_out[59],la_data_out[58],la_data_out[57],la_data_out[56],la_data_out[55],la_data_out[54],la_data_out[53],la_data_out[52],la_data_out[51],la_data_out[50],la_data_out[49],la_data_out[48],la_data_out[47],la_data_out[46],la_data_out[45],la_data_out[44],la_data_out[43],la_data_out[42],la_data_out[41],la_data_out[40],la_data_out[39],la_data_out[38],la_data_out[37],la_data_out[36],la_data_out[35],la_data_out[34],la_data_out[33],la_data_out[32],la_data_out[31],la_data_out[30],la_data_out[29],la_data_out[28],la_data_out[27],la_data_out[26],la_data_out[25],la_data_out[24],la_data_out[23],la_data_out[22],la_data_out[21],la_data_out[20],la_data_out[19],la_data_out[18],la_data_out[17],la_data_out[16],la_data_out[15],la_data_out[14],la_data_out[13],la_data_out[12],la_data_out[11],la_data_out[10],la_data_out[9],la_data_out[8],la_data_out[7],la_data_out[6],la_data_out[5],la_data_out[4],la_data_out[3],la_data_out[2],la_data_out[1],la_data_out[0]
*+ io_in[26],io_in[25],io_in[24],io_in[23],io_in[22],io_in[21],io_in[20],io_in[19],io_in[18],io_in[17],io_in[16],io_in[15],io_in[14],io_in[13],io_in[12],io_in[11],io_in[10],io_in[9],io_in[8],io_in[7],io_in[6],io_in[5],io_in[4],io_in[3],io_in[2],io_in[1],io_in[0]
*+ io_in_3v3[26],io_in_3v3[25],io_in_3v3[24],io_in_3v3[23],io_in_3v3[22],io_in_3v3[21],io_in_3v3[20],io_in_3v3[19],io_in_3v3[18],io_in_3v3[17],io_in_3v3[16],io_in_3v3[15],io_in_3v3[14],io_in_3v3[13],io_in_3v3[12],io_in_3v3[11],io_in_3v3[10],io_in_3v3[9],io_in_3v3[8],io_in_3v3[7],io_in_3v3[6],io_in_3v3[5],io_in_3v3[4],io_in_3v3[3],io_in_3v3[2],io_in_3v3[1],io_in_3v3[0] user_clock2
*+ io_out[26],io_out[25],io_out[24],io_out[23],io_out[22],io_out[21],io_out[20],io_out[19],io_out[18],io_out[17],io_out[16],io_out[15],io_out[14],io_out[13],io_out[12],io_out[11],io_out[10],io_out[9],io_out[8],io_out[7],io_out[6],io_out[5],io_out[4],io_out[3],io_out[2],io_out[1],io_out[0]
*+ io_oeb[26],io_oeb[25],io_oeb[24],io_oeb[23],io_oeb[22],io_oeb[21],io_oeb[20],io_oeb[19],io_oeb[18],io_oeb[17],io_oeb[16],io_oeb[15],io_oeb[14],io_oeb[13],io_oeb[12],io_oeb[11],io_oeb[10],io_oeb[9],io_oeb[8],io_oeb[7],io_oeb[6],io_oeb[5],io_oeb[4],io_oeb[3],io_oeb[2],io_oeb[1],io_oeb[0]
*+ gpio_analog[17],gpio_analog[16],gpio_analog[15],gpio_analog[14],gpio_analog[13],gpio_analog[12],gpio_analog[11],gpio_analog[10],gpio_analog[9],gpio_analog[8],gpio_analog[7],gpio_analog[6],gpio_analog[5],gpio_analog[4],gpio_analog[3],gpio_analog[2],gpio_analog[1],gpio_analog[0]
*+ gpio_noesd[17],gpio_noesd[16],gpio_noesd[15],gpio_noesd[14],gpio_noesd[13],gpio_noesd[12],gpio_noesd[11],gpio_noesd[10],gpio_noesd[9],gpio_noesd[8],gpio_noesd[7],gpio_noesd[6],gpio_noesd[5],gpio_noesd[4],gpio_noesd[3],gpio_noesd[2],gpio_noesd[1],gpio_noesd[0]
*+ io_analog[10],io_analog[9],io_analog[8],io_analog[7],io_analog[6],io_analog[5],io_analog[4],io_analog[3],io_analog[2],io_analog[1],io_analog[0] io_clamp_high[2],io_clamp_high[1],io_clamp_high[0] io_clamp_low[2],io_clamp_low[1],io_clamp_low[0]
*+ user_irq[2],user_irq[1],user_irq[0]
*+ la_oenb[127],la_oenb[126],la_oenb[125],la_oenb[124],la_oenb[123],la_oenb[122],la_oenb[121],la_oenb[120],la_oenb[119],la_oenb[118],la_oenb[117],la_oenb[116],la_oenb[115],la_oenb[114],la_oenb[113],la_oenb[112],la_oenb[111],la_oenb[110],la_oenb[109],la_oenb[108],la_oenb[107],la_oenb[106],la_oenb[105],la_oenb[104],la_oenb[103],la_oenb[102],la_oenb[101],la_oenb[100],la_oenb[99],la_oenb[98],la_oenb[97],la_oenb[96],la_oenb[95],la_oenb[94],la_oenb[93],la_oenb[92],la_oenb[91],la_oenb[90],la_oenb[89],la_oenb[88],la_oenb[87],la_oenb[86],la_oenb[85],la_oenb[84],la_oenb[83],la_oenb[82],la_oenb[81],la_oenb[80],la_oenb[79],la_oenb[78],la_oenb[77],la_oenb[76],la_oenb[75],la_oenb[74],la_oenb[73],la_oenb[72],la_oenb[71],la_oenb[70],la_oenb[69],la_oenb[68],la_oenb[67],la_oenb[66],la_oenb[65],la_oenb[64],la_oenb[63],la_oenb[62],la_oenb[61],la_oenb[60],la_oenb[59],la_oenb[58],la_oenb[57],la_oenb[56],la_oenb[55],la_oenb[54],la_oenb[53],la_oenb[52],la_oenb[51],la_oenb[50],la_oenb[49],la_oenb[48],la_oenb[47],la_oenb[46],la_oenb[45],la_oenb[44],la_oenb[43],la_oenb[42],la_oenb[41],la_oenb[40],la_oenb[39],la_oenb[38],la_oenb[37],la_oenb[36],la_oenb[35],la_oenb[34],la_oenb[33],la_oenb[32],la_oenb[31],la_oenb[30],la_oenb[29],la_oenb[28],la_oenb[27],la_oenb[26],la_oenb[25],la_oenb[24],la_oenb[23],la_oenb[22],la_oenb[21],la_oenb[20],la_oenb[19],la_oenb[18],la_oenb[17],la_oenb[16],la_oenb[15],la_oenb[14],la_oenb[13],la_oenb[12],la_oenb[11],la_oenb[10],la_oenb[9],la_oenb[8],la_oenb[7],la_oenb[6],la_oenb[5],la_oenb[4],la_oenb[3],la_oenb[2],la_oenb[1],la_oenb[0]
*.iopin vdda1
*.iopin vdda2
*.iopin vssa1
*.iopin vssa2
*.iopin vccd1
*.iopin vccd2
*.iopin vssd1
*.iopin vssd2
*.ipin wb_clk_i
*.ipin wb_rst_i
*.ipin wbs_stb_i
*.ipin wbs_cyc_i
*.ipin wbs_we_i
*.ipin wbs_sel_i[3],wbs_sel_i[2],wbs_sel_i[1],wbs_sel_i[0]
*.ipin
*+ wbs_dat_i[31],wbs_dat_i[30],wbs_dat_i[29],wbs_dat_i[28],wbs_dat_i[27],wbs_dat_i[26],wbs_dat_i[25],wbs_dat_i[24],wbs_dat_i[23],wbs_dat_i[22],wbs_dat_i[21],wbs_dat_i[20],wbs_dat_i[19],wbs_dat_i[18],wbs_dat_i[17],wbs_dat_i[16],wbs_dat_i[15],wbs_dat_i[14],wbs_dat_i[13],wbs_dat_i[12],wbs_dat_i[11],wbs_dat_i[10],wbs_dat_i[9],wbs_dat_i[8],wbs_dat_i[7],wbs_dat_i[6],wbs_dat_i[5],wbs_dat_i[4],wbs_dat_i[3],wbs_dat_i[2],wbs_dat_i[1],wbs_dat_i[0]
*.ipin
*+ wbs_adr_i[31],wbs_adr_i[30],wbs_adr_i[29],wbs_adr_i[28],wbs_adr_i[27],wbs_adr_i[26],wbs_adr_i[25],wbs_adr_i[24],wbs_adr_i[23],wbs_adr_i[22],wbs_adr_i[21],wbs_adr_i[20],wbs_adr_i[19],wbs_adr_i[18],wbs_adr_i[17],wbs_adr_i[16],wbs_adr_i[15],wbs_adr_i[14],wbs_adr_i[13],wbs_adr_i[12],wbs_adr_i[11],wbs_adr_i[10],wbs_adr_i[9],wbs_adr_i[8],wbs_adr_i[7],wbs_adr_i[6],wbs_adr_i[5],wbs_adr_i[4],wbs_adr_i[3],wbs_adr_i[2],wbs_adr_i[1],wbs_adr_i[0]
*.opin wbs_ack_o
*.opin
*+ wbs_dat_o[31],wbs_dat_o[30],wbs_dat_o[29],wbs_dat_o[28],wbs_dat_o[27],wbs_dat_o[26],wbs_dat_o[25],wbs_dat_o[24],wbs_dat_o[23],wbs_dat_o[22],wbs_dat_o[21],wbs_dat_o[20],wbs_dat_o[19],wbs_dat_o[18],wbs_dat_o[17],wbs_dat_o[16],wbs_dat_o[15],wbs_dat_o[14],wbs_dat_o[13],wbs_dat_o[12],wbs_dat_o[11],wbs_dat_o[10],wbs_dat_o[9],wbs_dat_o[8],wbs_dat_o[7],wbs_dat_o[6],wbs_dat_o[5],wbs_dat_o[4],wbs_dat_o[3],wbs_dat_o[2],wbs_dat_o[1],wbs_dat_o[0]
*.ipin
*+ la_data_in[127],la_data_in[126],la_data_in[125],la_data_in[124],la_data_in[123],la_data_in[122],la_data_in[121],la_data_in[120],la_data_in[119],la_data_in[118],la_data_in[117],la_data_in[116],la_data_in[115],la_data_in[114],la_data_in[113],la_data_in[112],la_data_in[111],la_data_in[110],la_data_in[109],la_data_in[108],la_data_in[107],la_data_in[106],la_data_in[105],la_data_in[104],la_data_in[103],la_data_in[102],la_data_in[101],la_data_in[100],la_data_in[99],la_data_in[98],la_data_in[97],la_data_in[96],la_data_in[95],la_data_in[94],la_data_in[93],la_data_in[92],la_data_in[91],la_data_in[90],la_data_in[89],la_data_in[88],la_data_in[87],la_data_in[86],la_data_in[85],la_data_in[84],la_data_in[83],la_data_in[82],la_data_in[81],la_data_in[80],la_data_in[79],la_data_in[78],la_data_in[77],la_data_in[76],la_data_in[75],la_data_in[74],la_data_in[73],la_data_in[72],la_data_in[71],la_data_in[70],la_data_in[69],la_data_in[68],la_data_in[67],la_data_in[66],la_data_in[65],la_data_in[64],la_data_in[63],la_data_in[62],la_data_in[61],la_data_in[60],la_data_in[59],la_data_in[58],la_data_in[57],la_data_in[56],la_data_in[55],la_data_in[54],la_data_in[53],la_data_in[52],la_data_in[51],la_data_in[50],la_data_in[49],la_data_in[48],la_data_in[47],la_data_in[46],la_data_in[45],la_data_in[44],la_data_in[43],la_data_in[42],la_data_in[41],la_data_in[40],la_data_in[39],la_data_in[38],la_data_in[37],la_data_in[36],la_data_in[35],la_data_in[34],la_data_in[33],la_data_in[32],la_data_in[31],la_data_in[30],la_data_in[29],la_data_in[28],la_data_in[27],la_data_in[26],la_data_in[25],la_data_in[24],la_data_in[23],la_data_in[22],la_data_in[21],la_data_in[20],la_data_in[19],la_data_in[18],la_data_in[17],la_data_in[16],la_data_in[15],la_data_in[14],la_data_in[13],la_data_in[12],la_data_in[11],la_data_in[10],la_data_in[9],la_data_in[8],la_data_in[7],la_data_in[6],la_data_in[5],la_data_in[4],la_data_in[3],la_data_in[2],la_data_in[1],la_data_in[0]
*.opin
*+ la_data_out[127],la_data_out[126],la_data_out[125],la_data_out[124],la_data_out[123],la_data_out[122],la_data_out[121],la_data_out[120],la_data_out[119],la_data_out[118],la_data_out[117],la_data_out[116],la_data_out[115],la_data_out[114],la_data_out[113],la_data_out[112],la_data_out[111],la_data_out[110],la_data_out[109],la_data_out[108],la_data_out[107],la_data_out[106],la_data_out[105],la_data_out[104],la_data_out[103],la_data_out[102],la_data_out[101],la_data_out[100],la_data_out[99],la_data_out[98],la_data_out[97],la_data_out[96],la_data_out[95],la_data_out[94],la_data_out[93],la_data_out[92],la_data_out[91],la_data_out[90],la_data_out[89],la_data_out[88],la_data_out[87],la_data_out[86],la_data_out[85],la_data_out[84],la_data_out[83],la_data_out[82],la_data_out[81],la_data_out[80],la_data_out[79],la_data_out[78],la_data_out[77],la_data_out[76],la_data_out[75],la_data_out[74],la_data_out[73],la_data_out[72],la_data_out[71],la_data_out[70],la_data_out[69],la_data_out[68],la_data_out[67],la_data_out[66],la_data_out[65],la_data_out[64],la_data_out[63],la_data_out[62],la_data_out[61],la_data_out[60],la_data_out[59],la_data_out[58],la_data_out[57],la_data_out[56],la_data_out[55],la_data_out[54],la_data_out[53],la_data_out[52],la_data_out[51],la_data_out[50],la_data_out[49],la_data_out[48],la_data_out[47],la_data_out[46],la_data_out[45],la_data_out[44],la_data_out[43],la_data_out[42],la_data_out[41],la_data_out[40],la_data_out[39],la_data_out[38],la_data_out[37],la_data_out[36],la_data_out[35],la_data_out[34],la_data_out[33],la_data_out[32],la_data_out[31],la_data_out[30],la_data_out[29],la_data_out[28],la_data_out[27],la_data_out[26],la_data_out[25],la_data_out[24],la_data_out[23],la_data_out[22],la_data_out[21],la_data_out[20],la_data_out[19],la_data_out[18],la_data_out[17],la_data_out[16],la_data_out[15],la_data_out[14],la_data_out[13],la_data_out[12],la_data_out[11],la_data_out[10],la_data_out[9],la_data_out[8],la_data_out[7],la_data_out[6],la_data_out[5],la_data_out[4],la_data_out[3],la_data_out[2],la_data_out[1],la_data_out[0]
*.ipin
*+ io_in[26],io_in[25],io_in[24],io_in[23],io_in[22],io_in[21],io_in[20],io_in[19],io_in[18],io_in[17],io_in[16],io_in[15],io_in[14],io_in[13],io_in[12],io_in[11],io_in[10],io_in[9],io_in[8],io_in[7],io_in[6],io_in[5],io_in[4],io_in[3],io_in[2],io_in[1],io_in[0]
*.ipin
*+ io_in_3v3[26],io_in_3v3[25],io_in_3v3[24],io_in_3v3[23],io_in_3v3[22],io_in_3v3[21],io_in_3v3[20],io_in_3v3[19],io_in_3v3[18],io_in_3v3[17],io_in_3v3[16],io_in_3v3[15],io_in_3v3[14],io_in_3v3[13],io_in_3v3[12],io_in_3v3[11],io_in_3v3[10],io_in_3v3[9],io_in_3v3[8],io_in_3v3[7],io_in_3v3[6],io_in_3v3[5],io_in_3v3[4],io_in_3v3[3],io_in_3v3[2],io_in_3v3[1],io_in_3v3[0]
*.ipin user_clock2
*.opin
*+ io_out[26],io_out[25],io_out[24],io_out[23],io_out[22],io_out[21],io_out[20],io_out[19],io_out[18],io_out[17],io_out[16],io_out[15],io_out[14],io_out[13],io_out[12],io_out[11],io_out[10],io_out[9],io_out[8],io_out[7],io_out[6],io_out[5],io_out[4],io_out[3],io_out[2],io_out[1],io_out[0]
*.opin
*+ io_oeb[26],io_oeb[25],io_oeb[24],io_oeb[23],io_oeb[22],io_oeb[21],io_oeb[20],io_oeb[19],io_oeb[18],io_oeb[17],io_oeb[16],io_oeb[15],io_oeb[14],io_oeb[13],io_oeb[12],io_oeb[11],io_oeb[10],io_oeb[9],io_oeb[8],io_oeb[7],io_oeb[6],io_oeb[5],io_oeb[4],io_oeb[3],io_oeb[2],io_oeb[1],io_oeb[0]
*.iopin
*+ gpio_analog[17],gpio_analog[16],gpio_analog[15],gpio_analog[14],gpio_analog[13],gpio_analog[12],gpio_analog[11],gpio_analog[10],gpio_analog[9],gpio_analog[8],gpio_analog[7],gpio_analog[6],gpio_analog[5],gpio_analog[4],gpio_analog[3],gpio_analog[2],gpio_analog[1],gpio_analog[0]
*.iopin
*+ gpio_noesd[17],gpio_noesd[16],gpio_noesd[15],gpio_noesd[14],gpio_noesd[13],gpio_noesd[12],gpio_noesd[11],gpio_noesd[10],gpio_noesd[9],gpio_noesd[8],gpio_noesd[7],gpio_noesd[6],gpio_noesd[5],gpio_noesd[4],gpio_noesd[3],gpio_noesd[2],gpio_noesd[1],gpio_noesd[0]
*.iopin
*+ io_analog[10],io_analog[9],io_analog[8],io_analog[7],io_analog[6],io_analog[5],io_analog[4],io_analog[3],io_analog[2],io_analog[1],io_analog[0]
*.iopin io_clamp_high[2],io_clamp_high[1],io_clamp_high[0]
*.iopin io_clamp_low[2],io_clamp_low[1],io_clamp_low[0]
*.opin user_irq[2],user_irq[1],user_irq[0]
*.ipin
*+ la_oenb[127],la_oenb[126],la_oenb[125],la_oenb[124],la_oenb[123],la_oenb[122],la_oenb[121],la_oenb[120],la_oenb[119],la_oenb[118],la_oenb[117],la_oenb[116],la_oenb[115],la_oenb[114],la_oenb[113],la_oenb[112],la_oenb[111],la_oenb[110],la_oenb[109],la_oenb[108],la_oenb[107],la_oenb[106],la_oenb[105],la_oenb[104],la_oenb[103],la_oenb[102],la_oenb[101],la_oenb[100],la_oenb[99],la_oenb[98],la_oenb[97],la_oenb[96],la_oenb[95],la_oenb[94],la_oenb[93],la_oenb[92],la_oenb[91],la_oenb[90],la_oenb[89],la_oenb[88],la_oenb[87],la_oenb[86],la_oenb[85],la_oenb[84],la_oenb[83],la_oenb[82],la_oenb[81],la_oenb[80],la_oenb[79],la_oenb[78],la_oenb[77],la_oenb[76],la_oenb[75],la_oenb[74],la_oenb[73],la_oenb[72],la_oenb[71],la_oenb[70],la_oenb[69],la_oenb[68],la_oenb[67],la_oenb[66],la_oenb[65],la_oenb[64],la_oenb[63],la_oenb[62],la_oenb[61],la_oenb[60],la_oenb[59],la_oenb[58],la_oenb[57],la_oenb[56],la_oenb[55],la_oenb[54],la_oenb[53],la_oenb[52],la_oenb[51],la_oenb[50],la_oenb[49],la_oenb[48],la_oenb[47],la_oenb[46],la_oenb[45],la_oenb[44],la_oenb[43],la_oenb[42],la_oenb[41],la_oenb[40],la_oenb[39],la_oenb[38],la_oenb[37],la_oenb[36],la_oenb[35],la_oenb[34],la_oenb[33],la_oenb[32],la_oenb[31],la_oenb[30],la_oenb[29],la_oenb[28],la_oenb[27],la_oenb[26],la_oenb[25],la_oenb[24],la_oenb[23],la_oenb[22],la_oenb[21],la_oenb[20],la_oenb[19],la_oenb[18],la_oenb[17],la_oenb[16],la_oenb[15],la_oenb[14],la_oenb[13],la_oenb[12],la_oenb[11],la_oenb[10],la_oenb[9],la_oenb[8],la_oenb[7],la_oenb[6],la_oenb[5],la_oenb[4],la_oenb[3],la_oenb[2],la_oenb[1],la_oenb[0]
x1 iref_cp2 vssa1 vdda1 net13 net12 net6 net1 net5 io_analog[10] io_analog[9] net4 net7 net2
+ gpio_noesd[7] net11 net14 net8 net9 net3 net10 net20 net15 net27 net21 net23 net25 net24 net18 net19 net22 net17
+ net26 net16 net28 top_pll_v1
x2 vdda1 io_analog[5] iref_cp0 iref_cp1 iref_cp2 net29 net30 iref4 iref2 iref3 iref1 iref0 bias
x3 iref_cp1 vssa1 vdda1 net43 net42 net36 net31 net35 io_analog[10] io_analog[8] net34 net37 net32
+ gpio_noesd[7] net41 net44 net38 net39 net33 net40 net50 net45 net57 net51 net53 net55 net54 net48 net49 net52
+ net47 net56 net46 net58 gpio_noesd[8] top_pll_v2
XC1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=9 m=9
XC2 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=9 m=9
XC3 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=7 m=7
XC4 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=15 m=15
XC5 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=15 m=15
XC6 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=15 m=15
XC7 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=15 m=15
XC8 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=15 m=15
XC9 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=15 m=15
x5 vdda1 io_analog[3] io_analog[2] io_analog[0] io_analog[1] vssa1 io_analog[6] gpio_noesd[4]
+ gpio_noesd[5] gpio_noesd[6] gpio_noesd[3] gpio_noesd[1] gpio_noesd[2] iref0 io_analog[4] iref1 iref2 iref3 iref4
+ res_amp_top
XC10 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=10 m=10
x4 iref_cp0 vssa1 vdda1 net71 net70 net64 net60 net92 io_analog[10] net63 io_analog[7] net62 net65
+ net59 gpio_noesd[7] net69 net72 net66 net67 net68 net61 gpio_noesd[10] gpio_noesd[11] gpio_noesd[9] net78
+ net73 net91 net79 net75 net74 net76 net77 net81 net90 net89 net88 net87 net86 net85 net84 net83 net82
+ net80 gpio_noesd[8] top_pll_v3
**.ends

* expanding   symbol:  top_pll_v1.sym # of pins=34
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/top_pll_v1.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/top_pll_v1.sch
.subckt top_pll_v1  iref_cp vss vdd vco_out vco_vctrl Up pfd_QA nUp in_ref out_to_pad Down nDown
+ pfd_QB vco_D0 lf_vc out_first_buffer cp_biasp cp_pswitch pfd_reset cp_nswitch out_by_2 out_to_div
+ out_div_by_5 n_out_by_2 div_5_nQ0 div_5_Q1_shift div_5_Q1 n_out_buffer_div_2 out_buffer_div_2 div_5_Q0
+ n_out_div_2 div_5_nQ2 out_div_2 out_to_buffer
*.iopin vdd
*.iopin vss
*.ipin in_ref
*.iopin pfd_QA
*.iopin pfd_QB
*.iopin Up
*.iopin nUp
*.iopin Down
*.iopin nDown
*.iopin pfd_reset
*.iopin cp_nswitch
*.iopin cp_pswitch
*.iopin cp_biasp
*.ipin iref_cp
*.iopin lf_vc
*.iopin vco_D0
*.iopin vco_vctrl
*.iopin vco_out
*.iopin out_first_buffer
*.iopin out_to_buffer
*.iopin out_to_div
*.iopin out_by_2
*.iopin n_out_by_2
*.iopin out_div_2
*.iopin n_out_div_2
*.iopin out_buffer_div_2
*.iopin n_out_buffer_div_2
*.iopin div_5_Q1
*.iopin div_5_Q1_shift
*.iopin div_5_nQ0
*.iopin div_5_Q0
*.iopin div_5_nQ2
*.iopin out_div_by_5
*.iopin out_to_pad
x1 vss vdd pfd_QA in_ref out_div_by_5 pfd_QB pfd_reset PFD
x2 vdd Up nUp vco_vctrl Down nDown vss iref_cp cp_nswitch cp_pswitch cp_biasp charge_pump
x3 Up vdd pfd_QA nUp Down pfd_QB vss nDown pfd_cp_interface
x4 vss vco_vctrl lf_vc loop_filter
x5 vdd vco_out vco_D0 vco_vctrl vss csvco
x6 vdd vco_out out_to_buffer out_to_div vss out_first_buffer ring_osc_buffer
x7 vdd out_div_by_5 out_by_2 vss n_out_by_2 div_5_nQ2 div_5_Q1 div_5_nQ0 div_5_Q0 div_5_Q1_shift
+ div_by_5
x8 n_out_by_2 vss out_to_div vdd out_by_2 out_div_2 n_out_div_2 out_buffer_div_2 n_out_buffer_div_2
+ div_by_2
x9 vdd out_to_pad out_to_buffer vss buffer_salida
.ends


* expanding   symbol:  bias.sym # of pins=12
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/bias.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/bias.sch
.subckt bias  vdd iref iref_0 iref_1 iref_2 iref_3 iref_4 iref_5 iref_6 iref_7 iref_8 iref_9
*.iopin iref
*.iopin vdd
*.opin iref_0
*.opin iref_1
*.opin iref_2
*.opin iref_3
*.opin iref_4
*.opin iref_5
*.opin iref_6
*.opin iref_7
*.opin iref_8
*.opin iref_9
XM1 iref iref vbp1 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM2 vbp1 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM3 net1 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM4 iref_0 iref net1 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM5 net2 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM6 iref_1 iref net2 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM7 net3 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM8 iref_2 iref net3 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM9 net4 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM10 iref_3 iref net4 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM11 net5 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM12 iref_4 iref net5 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM13 net6 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM14 iref_5 iref net6 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM15 net7 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM16 iref_6 iref net7 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM17 net8 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM18 iref_7 iref net8 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM19 net9 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM20 iref_8 iref net9 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM21 net10 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
XM22 iref_9 iref net10 vdd sky130_fd_pr__pfet_01v8_lvt L=0.45 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=25 m=25 
.ends


* expanding   symbol:  top_pll_v2.sym # of pins=35
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/top_pll_v2.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/top_pll_v2.sch
.subckt top_pll_v2  iref_cp vss vdd vco_out vco_vctrl Up pfd_QA nUp in_ref out_to_pad Down nDown
+ pfd_QB D0_vco lf_vc out_first_buffer cp_biasp cp_pswitch pfd_reset cp_nswitch out_by_2 out_to_div
+ out_div_by_5 n_out_by_2 div_5_nQ0 div_5_Q1_shift div_5_Q1 n_out_buffer_div_2 out_buffer_div_2 div_5_Q0
+ n_out_div_2 div_5_nQ2 out_div_2 out_to_buffer D0_cap
*.iopin vdd
*.iopin vss
*.ipin in_ref
*.iopin pfd_QA
*.iopin pfd_QB
*.iopin Up
*.iopin nUp
*.iopin Down
*.iopin nDown
*.iopin pfd_reset
*.iopin cp_nswitch
*.iopin cp_pswitch
*.iopin cp_biasp
*.ipin iref_cp
*.iopin lf_vc
*.iopin D0_vco
*.iopin vco_vctrl
*.iopin vco_out
*.iopin out_first_buffer
*.iopin out_to_buffer
*.iopin out_to_div
*.iopin out_by_2
*.iopin n_out_by_2
*.iopin out_div_2
*.iopin n_out_div_2
*.iopin out_buffer_div_2
*.iopin n_out_buffer_div_2
*.iopin div_5_Q1
*.iopin div_5_Q1_shift
*.iopin div_5_nQ0
*.iopin div_5_Q0
*.iopin div_5_nQ2
*.iopin out_div_by_5
*.iopin out_to_pad
*.ipin D0_cap
x1 vss vdd pfd_QA in_ref out_div_by_5 pfd_QB pfd_reset PFD
x2 vdd Up nUp vco_vctrl Down nDown vss iref_cp cp_nswitch cp_pswitch cp_biasp charge_pump
x3 Up vdd pfd_QA nUp Down pfd_QB vss nDown pfd_cp_interface
x5 vdd vco_out D0_vco vco_vctrl vss csvco
x6 vdd vco_out out_to_buffer out_to_div vss out_first_buffer ring_osc_buffer
x7 vdd out_div_by_5 out_by_2 vss n_out_by_2 div_5_nQ2 div_5_Q1 div_5_nQ0 div_5_Q0 div_5_Q1_shift
+ div_by_5
x8 n_out_by_2 vss out_to_div vdd out_by_2 out_div_2 n_out_div_2 out_buffer_div_2 n_out_buffer_div_2
+ div_by_2
x9 vdd out_to_pad out_to_buffer vss buffer_salida
x4 vss vco_vctrl lf_vc D0_cap loop_filter_v2
.ends


* expanding   symbol:  res_amp_top.sym # of pins=19
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/res_amp_top.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/res_amp_top.sch
.subckt res_amp_top  avdd1p8 inp inn outp outn avss1p8 clkp iref_reg0 iref_reg1 iref_reg2 delay_reg0
+ delay_reg2 delay_reg1 iref0 clkn iref1 iref2 iref3 iref4
*.ipin inp
*.ipin inn
*.ipin clkp
*.ipin clkn
*.iopin avdd1p8
*.iopin avss1p8
*.ipin iref0
*.ipin iref1
*.ipin iref2
*.ipin iref3
*.ipin iref4
*.opin outn
*.opin outp
*.ipin iref_reg0
*.ipin iref_reg1
*.ipin iref_reg2
*.ipin delay_reg0
*.ipin delay_reg1
*.ipin delay_reg2
x2 avdd1p8 rst inp inn outp_amp outn_amp avss1p8 outp_cap outn_cap clk_amp iref_reg0 iref_reg1
+ iref_reg2 delay_reg0 delay_reg2 delay_reg1 iref0 res_amp_lin_prog
x1 avdd1p8 clkp clkn avss1p8 clk_amp rst res_amp_sync_v2
x3 avdd1p8 iref1 outp_cap outp avss1p8 outn_cap outn iref2 iref3 iref4 source_follower_buff_diff
XC1 outp_cap avss1p8 sky130_fd_pr__cap_mim_m3_1 W=5.5 L=7.5 MF=1 m=1
XC2 outn_cap avss1p8 sky130_fd_pr__cap_mim_m3_1 W=5.5 L=7.5 MF=1 m=1
.ends


* expanding   symbol:  top_pll_v3.sym # of pins=44
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/top_pll_v3.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/top_pll_v3.sch
.subckt top_pll_v3  iref_cp vss vdd vco_out vco_vctrl Up pfd_QA out_to_buffer in_ref nUp out_to_pad
+ Down nDown pfd_QB vco_D0 lf_vc out_first_buffer cp_biasp cp_pswitch cp_nswitch pfd_reset s_0 MC s_1
+ out_by_2 out_to_div out_div n_out_by_2 n_out_div_2 out_div_2 n_out_buffer_div_2 out_buffer_div_2 n_clk_0 s1n
+ s0n clk_2_f clk_d clk_out_mux21 clk_5 clk_pre n_clk_1 clk_1 clk_0 lf_D0
*.iopin vdd
*.iopin vss
*.ipin in_ref
*.iopin pfd_QA
*.iopin pfd_QB
*.iopin Up
*.iopin nUp
*.iopin Down
*.iopin nDown
*.iopin pfd_reset
*.iopin cp_nswitch
*.iopin cp_pswitch
*.iopin cp_biasp
*.ipin iref_cp
*.iopin lf_vc
*.ipin vco_D0
*.iopin vco_vctrl
*.iopin vco_out
*.iopin out_first_buffer
*.iopin out_to_buffer
*.iopin out_to_div
*.iopin out_by_2
*.iopin n_out_by_2
*.iopin out_div_2
*.iopin n_out_div_2
*.iopin out_buffer_div_2
*.iopin n_out_buffer_div_2
*.iopin out_div
*.opin out_to_pad
*.iopin clk_0
*.iopin n_clk_0
*.iopin clk_1
*.iopin n_clk_1
*.iopin clk_pre
*.iopin clk_5
*.iopin clk_out_mux21
*.iopin clk_d
*.iopin clk_2_f
*.iopin s0n
*.iopin s1n
*.ipin MC
*.ipin s_0
*.ipin s_1
*.ipin lf_D0
x1 vss vdd pfd_QA in_ref out_div pfd_QB pfd_reset PFD
x2 Up vdd pfd_QA nUp Down pfd_QB vss nDown pfd_cp_interface
x3 vdd Up nUp vco_vctrl Down nDown vss iref_cp cp_nswitch cp_pswitch cp_biasp charge_pump
x5 vdd vco_out vco_D0 vco_vctrl vss csvco
x6 vdd vco_out out_to_buffer out_to_div vss out_first_buffer ring_osc_buffer
x7 vdd out_to_pad out_to_buffer vss buffer_salida
x8 n_out_by_2 vss out_to_div vdd out_by_2 out_div_2 n_out_div_2 out_buffer_div_2 n_out_buffer_div_2
+ div_by_2
x9 s1n s0n s_0 s_1 MC clk_0 clk_pre vss vdd clk_out_mux21 clk_d n_clk_0 out_div out_by_2 clk_5
+ clk_2_f n_out_by_2 clk_1 n_clk_1 freq_div
x4 vss vco_vctrl lf_vc lf_D0 loop_filter_v2
.ends


* expanding   symbol:  PFD.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/PFD.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/PFD.sch
.subckt PFD  vss vdd Up A B Down Reset
*.iopin vdd
*.iopin vss
*.ipin A
*.ipin B
*.opin Down
*.opin Up
*.iopin Reset
x1 vdd A Up Reset vss DFF
x2 vdd B Down Reset vss DFF
x3 vdd Reset Up Down vss and_pfd
.ends


* expanding   symbol:  charge_pump.sym # of pins=11
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/charge_pump.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/charge_pump.sch
.subckt charge_pump  vdd Up nUp out Down nDown vss iref nswitch pswitch biasp
*.iopin vss
*.iopin vdd
*.ipin Down
*.ipin nUp
*.ipin Up
*.ipin nDown
*.opin out
*.iopin nswitch
*.iopin pswitch
*.ipin iref
*.iopin biasp
XM1 out pswitch vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=25 m=25 
XM2 out nswitch vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=25 m=25 
XM3 pswitch nUp biasp vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10 
XM4 pswitch Up vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10 
XM5 nswitch Down iref vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10 
XM6 nswitch nDown vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10 
XM7 pswitch nUp pswitch vdd sky130_fd_pr__pfet_01v8 L=2 W=4.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10 
XM8 nswitch Down nswitch vss sky130_fd_pr__nfet_01v8 L=1.5 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10 
XM9 iref iref vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=25 m=25 
XM10 biasp iref vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=25 m=25 
XM11 biasp biasp vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=25 m=25 
.ends


* expanding   symbol:  pfd_cp_interface.sym # of pins=8
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/pfd_cp_interface.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/pfd_cp_interface.sch
.subckt pfd_cp_interface  Up vdd QA nUp Down QB vss nDown
*.iopin vdd
*.iopin vss
*.ipin QA
*.ipin QB
*.opin nDown
*.opin Down
*.opin nUp
*.opin Up
x5 vdd nDown nQB vss trans_gate
x3 vdd Up nQA vss inverter_cp_x1
x1 vdd nQB QB vss inverter_cp_x1
x2 vdd nQA QA vss inverter_cp_x1
x4 vdd nUp Up vss inverter_cp_x2
x6 vdd Down nDown vss inverter_cp_x2
.ends


* expanding   symbol:  loop_filter.sym # of pins=3
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/loop_filter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/loop_filter.sch
.subckt loop_filter  vss in vc_pex
*.iopin in
*.iopin vss
*.iopin vc_pex
x1 in net1 vss res_loop_filter
x2 vc_pex net1 vss res_loop_filter
x3 vc_pex net1 vss res_loop_filter
x4 vc_pex vss cap1_loop_filter
x5 in vss cap2_loop_filter
.ends


* expanding   symbol:  csvco.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/csvco.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/csvco.sch
.subckt csvco  vdd out D0 vctrl vss
*.ipin vctrl
*.iopin vss
*.iopin vdd
*.opin out
*.ipin D0
XM1 vbp vctrl vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 vbp vbp vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x1 vdd vbp out out1 vctrl vss D0 csvco_branch
x2 vdd vbp out1 out2 vctrl vss D0 csvco_branch
x3 vdd vbp out2 out vctrl vss D0 csvco_branch
.ends


* expanding   symbol:  ring_osc_buffer.sym # of pins=6
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/ring_osc_buffer.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/ring_osc_buffer.sch
.subckt ring_osc_buffer  vdd in_vco out_pad out_div vss o1
*.iopin vdd
*.iopin vss
*.ipin in_vco
*.opin out_pad
*.opin out_div
*.iopin o1
x1 vdd o1 in_vco vss inverter_min_x2
x2 vdd out_div o1 vss inverter_min_x4
x3 vdd out_pad out_div vss inverter_min_x4
.ends


* expanding   symbol:  div_by_5.sym # of pins=10
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/div_by_5.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/div_by_5.sch
.subckt div_by_5  vdd CLK_5 CLK vss nCLK nQ2 Q1 nQ0 Q0 Q1_shift
*.iopin vdd
*.iopin vss
*.ipin CLK
*.opin CLK_5
*.ipin nCLK
*.iopin nQ2
*.iopin Q1
*.iopin Q0
*.iopin nQ0
*.iopin Q1_shift
x8 Q1 Q0 vss vss vdd vdd D2 sky130_fd_sc_hs__and2_1
x9 Q1 Q0 vss vss vdd vdd D1 sky130_fd_sc_hs__xor2_1
x10 nQ2 nQ0 vss vss vdd vdd D0 sky130_fd_sc_hs__and2_1
x12 Q1 Q1_shift vss vss vdd vdd CLK_5 sky130_fd_sc_hs__or2_1
x1 vdd Q2 nQ2 vss D2 CLK nCLK DFlipFlop
x2 vdd Q1 nQ1 vss D1 CLK nCLK DFlipFlop
x3 vdd Q0 nQ0 vss D0 CLK nCLK DFlipFlop
x4 vdd Q1_shift nQ1_shift vss Q1 nCLK CLK DFlipFlop
.ends


* expanding   symbol:  div_by_2.sym # of pins=9
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/div_by_2.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/div_by_2.sch
.subckt div_by_2  nCLK_2 vss CLK vdd CLK_2 out_div nout_div o1 o2
*.ipin CLK
*.opin CLK_2
*.iopin vss
*.iopin vdd
*.opin nCLK_2
*.iopin nout_div
*.iopin o2
*.iopin o1
*.iopin out_div
x1 vdd out_div nout_div vss nout_div CLK_d nCLK_d DFlipFlop
x2 vdd CLK_d CLK nCLK_d vss clock_inverter
x3 vdd o1 out_div vss inverter_min_x2
x4 vdd CLK_2 o1 vss inverter_min_x4
x5 vdd o2 nout_div vss inverter_min_x2
x6 vdd nCLK_2 o2 vss inverter_min_x4
.ends


* expanding   symbol:  buffer_salida.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/buffer_salida.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/buffer_salida.sch
.subckt buffer_salida  vdd out in vss
*.iopin vss
*.ipin in
*.iopin vdd
*.opin out
XM2 net1 in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM1 net1 in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM3 net2 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=32 m=32 
XM4 net2 net1 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=32 m=32 
XM5 out net2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=256 m=256 
XM6 out net2 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=256 m=256 
.ends


* expanding   symbol:  loop_filter_v2.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/loop_filter_v2.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/loop_filter_v2.sch
.subckt loop_filter_v2  vss in vc_pex D0_cap
*.iopin in
*.iopin vss
*.iopin vc_pex
*.iopin D0_cap
x1 in net1 vss res_loop_filter
x2 vc_pex net1 vss res_loop_filter
x3 vc_pex net1 vss res_loop_filter
x4 vc_pex vss cap1_loop_filter
x5 in vss cap2_loop_filter
XM1 in D0_cap net2 vss sky130_fd_pr__nfet_01v8 L=0.3 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x6 net2 vss cap3_loop_filter
.ends


* expanding   symbol:  res_amp_lin_prog.sym # of pins=17
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/res_amp_lin_prog.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/res_amp_lin_prog.sch
.subckt res_amp_lin_prog  avdd1p8 rst inp inn outp outn avss1p8 outp_cap outn_cap clk iref_reg0
+ iref_reg1 iref_reg2 delay_reg0 delay_reg2 delay_reg1 iref
*.ipin clk
*.opin outp
*.opin outn
*.iopin avdd1p8
*.iopin avss1p8
*.ipin iref
*.ipin inp
*.ipin inn
*.ipin iref_reg0
*.ipin iref_reg1
*.ipin iref_reg2
*.opin outp_cap
*.opin outn_cap
*.ipin delay_reg0
*.ipin delay_reg1
*.ipin delay_reg2
*.ipin rst
x3 avdd1p8 clk avss1p8 clk_out delay_reg0 delay_reg1 delay_reg2 delay_cell_buff
XM3 outn_cap rst avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3 
x4 avdd1p8 clk_out inp inn outp outn avss1p8 vctrl res_amp_lin
XM1 outp clk_out_b outp_cap avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5 
XM2 outn clk_out_b outn_cap avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5 
XM5 outp_cap clk_out outp avdd1p8 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10 
XM6 outn_cap clk_out outn avdd1p8 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10 
x5 avdd1p8 clk_out_b clk_out avss1p8 inverter_min_x4
XM4 outp_cap rst avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3 
x7 avdd1p8 iref avss1p8 vctrl iref_reg0 iref_reg1 iref_reg2 iref_ctrl_res_amp
.ends


* expanding   symbol:  res_amp_sync_v2.sym # of pins=6
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/res_amp_sync_v2.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/res_amp_sync_v2.sch
.subckt res_amp_sync_v2  avdd1p8 clkp clkn avss1p8 clk_amp rst
*.ipin clkn
*.ipin clkp
*.iopin avdd1p8
*.iopin avss1p8
*.opin rst
*.opin clk_amp
x4 avdd1p8 net1 net3 net2 avss1p8 nand_logic
x1 avdd1p8 d1 q1 avss1p8 inverter_min_x4
x5 avdd1p8 pulse net3 avss1p8 inverter_min_x4
x21 avdd1p8 pulse net6 clkp avss1p8 nand_logic
x3 avdd1p8 net2 net7 avss1p8 d1 clkp clkn DFlipFlop
x6 avdd1p8 net1 net8 avss1p8 q2 clkp clkn DFlipFlop
x7 avdd1p8 q1 net9 avss1p8 d1 clkp clkn DFlipFlop
x8 avdd1p8 q2 net10 avss1p8 d2 d1 q1 DFlipFlop
x9 avdd1p8 net4 net11 avss1p8 pulse clkp clkn DFlipFlop
x2 avdd1p8 d2 q2 avss1p8 inverter_min_x4
x10 avdd1p8 rst net6 avss1p8 inverter_min_x4
x11 avdd1p8 net5 net4 avss1p8 inverter_min_x4
x12 avdd1p8 clk_amp net5 avss1p8 inverter_min_x16
.ends


* expanding   symbol:  source_follower_buff_diff.sym # of pins=10
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/source_follower_buff_diff.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/source_follower_buff_diff.sch
.subckt source_follower_buff_diff  avdd1p8 iref1 inp outp avss1p8 inn outn iref2 iref3 iref4
*.iopin avdd1p8
*.iopin avss1p8
*.opin outp
*.opin outn
*.ipin inp
*.ipin inn
*.ipin iref1
*.ipin iref2
*.ipin iref3
*.ipin iref4
x1 avdd1p8 iref1 inp outp_int avss1p8 source_follower_buff_pmos
x2 avdd1p8 iref2 outp_int outp avss1p8 source_follower_buff_nmos
x3 avdd1p8 iref3 inn outn_int avss1p8 source_follower_buff_pmos
x4 avdd1p8 iref4 outn_int outn avss1p8 source_follower_buff_nmos
.ends


* expanding   symbol:  freq_div.sym # of pins=19
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/freq_div.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/freq_div.sch
.subckt freq_div  s_1_n s_0_n s_0 s_1 MC clk_0 clk_pre vss vdd clk_out_mux21 clk_d n_clk_0 out in_a
+ clk_5 clk_2 in_b clk_1 n_clk_1
*.ipin s_0
*.iopin vdd
*.iopin vss
*.ipin in_a
*.ipin in_b
*.opin out
*.ipin MC
*.ipin s_1
*.iopin clk_0
*.iopin n_clk_0
*.iopin clk_1
*.iopin n_clk_1
*.iopin clk_pre
*.iopin clk_5
*.iopin clk_out_mux21
*.iopin clk_d
*.iopin clk_2
*.iopin s_0_n
*.iopin s_1_n
x2 vdd clk_pre clk_0 n_clk_0 vss MC net2 net1 net3 net4 prescaler_23
x3 net14 vss clk_out_mux21 vdd clk_2 net5 net6 net7 net8 div_by_2
x4 vdd clk_5 clk_1 vss n_clk_1 net9 net10 net12 net13 net11 div_by_5
x9 vdd s_0_n s_0 vss inverter_min_x2
x1 vdd vss in_a in_b n_clk_0 clk_0 s_0 n_clk_1 clk_1 s_0_n mux2to4
x6 vdd vss clk_out_mux21 clk_pre s_0 clk_5 s_0_n mux2to1
x5 vdd vss out clk_d s_1 clk_2 s_1_n mux2to1
x7 vdd s_1_n s_1 vss inverter_min_x2
x8 vdd net15 clk_out_mux21 vss inverter_min_x2
x10 vdd clk_d net15 vss inverter_min_x4
.ends


* expanding   symbol:  DFF.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/DFF.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/DFF.sch
.subckt DFF  D CLK Q Reset vss
*.ipin D
*.ipin CLK
*.opin Q
*.ipin Reset
*.iopin vss
x1 D CLK Q P vss nor
x2 D P P1 Q vss nor
x3 D P P2 P1 vss nor
x4 D P1 Reset P2 vss nor
.ends


* expanding   symbol:  and_pfd.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/and_pfd.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/and_pfd.sch
.subckt and_pfd  vdd out A B vss
*.iopin vdd
*.iopin vss
*.opin out
*.ipin A
*.ipin B
XM1 out_nand A net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out_nand A vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net1 B vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 out_nand B net2 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 net2 A vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 out_nand B vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 out out_nand vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 out out_nand vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  trans_gate.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/trans_gate.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/trans_gate.sch
.subckt trans_gate  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out vss in vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM1 out vdd in vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
.ends


* expanding   symbol:  inverter_cp_x1.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_cp_x1.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_cp_x1.sch
.subckt inverter_cp_x1  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
.ends


* expanding   symbol:  inverter_cp_x2.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_cp_x2.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_cp_x2.sch
.subckt inverter_cp_x2  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
.ends


* expanding   symbol:  res_loop_filter.sym # of pins=3
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/res_loop_filter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/res_loop_filter.sch
.subckt res_loop_filter  in out vss
*.iopin in
*.iopin vss
*.iopin out
XR3 out in vss sky130_fd_pr__res_high_po_5p73 L=22.92 mult=1 m=1
.ends


* expanding   symbol:  cap1_loop_filter.sym # of pins=2
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/cap1_loop_filter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/cap1_loop_filter.sch
.subckt cap1_loop_filter  in out
*.iopin in
*.iopin out
XC1 in out sky130_fd_pr__cap_mim_m3_1 W=25 L=25 MF=25 m=25
.ends


* expanding   symbol:  cap2_loop_filter.sym # of pins=2
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/cap2_loop_filter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/cap2_loop_filter.sch
.subckt cap2_loop_filter  in out
*.iopin in
*.iopin out
XC1 in out sky130_fd_pr__cap_mim_m3_1 W=20 L=20 MF=9 m=9
.ends


* expanding   symbol:  csvco_branch.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/csvco_branch.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/csvco_branch.sch
.subckt csvco_branch  vdd vbp in out vctrl vss D0
*.ipin vctrl
*.ipin vbp
*.iopin vdd
*.iopin vss
*.ipin in
*.opin out
*.ipin D0
XM1 vdd_inv vbp vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10 
XM2 vss_inv vctrl vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10 
XM4 out D0 net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x1 vdd_inv out in vss_inv vdd vss inverter_csvco
C1 net1 vss 5.78f m=1
.ends


* expanding   symbol:  inverter_min_x2.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_min_x2.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_min_x2.sch
.subckt inverter_min_x2  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:  inverter_min_x4.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_min_x4.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_min_x4.sch
.subckt inverter_min_x4  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
.ends


* expanding   symbol:  DFlipFlop.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/DFlipFlop.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/DFlipFlop.sch
.subckt DFlipFlop  vdd Q nQ vss D CLK nCLK
*.iopin vdd
*.iopin vss
*.opin Q
*.opin nQ
*.ipin D
*.ipin CLK
*.ipin nCLK
x1 vdd D_d D nD_d vss clock_inverter
x2 vdd nA A D_d nD_d CLK vss latch_diff
x3 vdd nQ Q A nA nCLK vss latch_diff
.ends


* expanding   symbol:  clock_inverter.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/clock_inverter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/clock_inverter.sch
.subckt clock_inverter  vdd CLK_d CLK nCLK_d vss
*.ipin CLK
*.iopin vdd
*.iopin vss
*.opin nCLK_d
*.opin CLK_d
x5 vdd nCLK_d net1 vss trans_gate
x1 vdd CLK_d net2 vss inverter_cp_x1
x2 vdd net2 CLK vss inverter_cp_x1
x3 vdd net1 CLK vss inverter_cp_x1
.ends


* expanding   symbol:  cap3_loop_filter.sym # of pins=2
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/cap3_loop_filter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/cap3_loop_filter.sch
.subckt cap3_loop_filter  in out
*.iopin in
*.iopin out
XC1 in out sky130_fd_pr__cap_mim_m3_1 W=20 L=20 MF=4 m=4
.ends


* expanding   symbol:  delay_cell_buff.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/delay_cell_buff.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/delay_cell_buff.sch
.subckt delay_cell_buff  avdd1p8 clk avss1p8 clk_out reg0 reg1 reg2
*.ipin clk
*.iopin avdd1p8
*.iopin avss1p8
*.opin clk_out
*.ipin reg2
*.ipin reg1
*.ipin reg0
x1 avdd1p8 reg2 avss1p8 clk3 net1 clk2 mux_2to1_logic
x2 avdd1p8 reg2 avss1p8 clk1 net2 clk mux_2to1_logic
x3 avdd1p8 reg1 avss1p8 net1 net3 net2 mux_2to1_logic
x4 avdd1p8 out_mux clk_out clk avss1p8 nand_logic
x513 avdd1p8 clk avss1p8 clk1_int buffer_no_inv_x05
x512 avdd1p8 clk1_int avss1p8 clk1 buffer_no_inv_x05
x511 avdd1p8 clk1 avss1p8 clk2_int buffer_no_inv_x05
x510 avdd1p8 clk2_int avss1p8 clk2 buffer_no_inv_x05
x59 avdd1p8 clk2 avss1p8 clk3_int buffer_no_inv_x05
x58 avdd1p8 clk3_int avss1p8 clk3 buffer_no_inv_x05
x57 avdd1p8 clk3 avss1p8 clk4_int buffer_no_inv_x05
x56 avdd1p8 clk4_int avss1p8 clk4 buffer_no_inv_x05
x55 avdd1p8 clk4 avss1p8 clk5_int buffer_no_inv_x05
x54 avdd1p8 clk5_int avss1p8 clk5 buffer_no_inv_x05
x53 avdd1p8 clk5 avss1p8 clk6_int buffer_no_inv_x05
x52 avdd1p8 clk6_int avss1p8 clk6 buffer_no_inv_x05
x51 avdd1p8 clk6 avss1p8 clk7_int buffer_no_inv_x05
x50 avdd1p8 clk7_int avss1p8 clk7 buffer_no_inv_x05
x5 avdd1p8 reg2 avss1p8 clk7 net4 clk6 mux_2to1_logic
x6 avdd1p8 reg2 avss1p8 clk5 net5 clk4 mux_2to1_logic
x7 avdd1p8 reg1 avss1p8 net4 net6 net5 mux_2to1_logic
x8 avdd1p8 reg0 avss1p8 net6 out_mux net3 mux_2to1_logic
.ends


* expanding   symbol:  res_amp_lin.sym # of pins=8
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/res_amp_lin.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/res_amp_lin.sch
.subckt res_amp_lin  avdd1p8 clk inp inn outp outn avss1p8 vctrl
*.iopin avdd1p8
*.iopin avss1p8
*.opin outp
*.opin outn
*.ipin inn
*.ipin inp
*.ipin clk
*.ipin vctrl
XM6 int clk avdd1p8 avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3 
XM8 outn clk avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM9 outp clk avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 vp vctrl int avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5 
XM1 outn inp vp avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM2 outp inn vp avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
.ends


* expanding   symbol:  iref_ctrl_res_amp.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/iref_ctrl_res_amp.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/iref_ctrl_res_amp.sch
.subckt iref_ctrl_res_amp  avdd1p8 iref avss1p8 vctrl reg0 reg1 reg2
*.iopin avdd1p8
*.iopin avss1p8
*.ipin reg0
*.ipin reg1
*.ipin reg2
*.opin vctrl
*.ipin iref
XM7 iref iref net1 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM8 vctrl iref net2 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3 
XM9 vctrl vctrl net3 avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM10 net3 avss1p8 avdd1p8 avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3 
XM1 vctrl iref net4 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM2 vctrl iref net5 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4 
XM3 net4 reg0 avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM4 net5 reg1 avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4 
XM5 net2 avdd1p8 avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3 
XM6 net1 avdd1p8 avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM11 vctrl iref net6 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XM12 net6 reg2 avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
.ends


* expanding   symbol:  nand_logic.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/nand_logic.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/nand_logic.sch
.subckt nand_logic  avdd1p8 in1 out in2 avss1p8
*.ipin in1
*.ipin in2
*.opin out
*.iopin avdd1p8
*.iopin avss1p8
XM4 out in2 avdd1p8 avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1.02 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM5 n1 in1 avss1p8 avss1p8 sky130_fd_pr__nfet_01v8 L=0.15 W=1.02 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM1 out in2 n1 avss1p8 sky130_fd_pr__nfet_01v8 L=0.15 W=1.02 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 out in1 avdd1p8 avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1.02 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:  inverter_min_x16.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_min_x16.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_min_x16.sch
.subckt inverter_min_x16  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
.ends


* expanding   symbol:  source_follower_buff_pmos.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/source_follower_buff_pmos.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/source_follower_buff_pmos.sch
.subckt source_follower_buff_pmos  avdd1p8 iref in out avss1p8
*.iopin avdd1p8
*.iopin avss1p8
*.opin out
*.ipin in
*.ipin iref
XM5 net1 net1 avdd1p8 avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=15 m=15 
XM6 out net1 avdd1p8 avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=15 m=15 
XM1 avss1p8 in out avdd1p8 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20 
XM2 iref iref avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM3 net1 iref avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
.ends


* expanding   symbol:  source_follower_buff_nmos.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/source_follower_buff_nmos.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/source_follower_buff_nmos.sch
.subckt source_follower_buff_nmos  avdd1p8 iref in out avss1p8
*.iopin avdd1p8
*.iopin avss1p8
*.opin out
*.ipin in
*.ipin iref
XM2 net1 iref avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM1 out iref avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=160 m=160 
XM3 avdd1p8 in out avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=80 m=80 
XM4 iref iref net1 avss1p8 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
.ends


* expanding   symbol:  prescaler_23.sym # of pins=10
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/prescaler_23.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/prescaler_23.sch
.subckt prescaler_23  vdd CLK_23 CLK nCLK vss MC Q1 nCLK_23 Q2 Q2_d
*.iopin vdd
*.ipin CLK
*.ipin nCLK
*.ipin MC
*.iopin vss
*.opin CLK_23
*.iopin nCLK_23
*.iopin Q1
*.iopin Q2
*.iopin Q2_d
x3 nCLK_23 1 vss vss vdd vdd 2 sky130_fd_sc_hs__and2_1
x4 Q1 MC vss vss vdd vdd 1 sky130_fd_sc_hs__or2_1
x6 3 nCLK_23 MC vss vss vdd vdd CLK_23 sky130_fd_sc_hs__mux2_1
x7 Q2 Q2_d vss vss vdd vdd 3 sky130_fd_sc_hs__or2_1
x1 vdd Q1 net1 vss nCLK_23 CLK nCLK DFlipFlop
x2 vdd Q2 nCLK_23 vss 2 CLK nCLK DFlipFlop
x5 vdd Q2_d net2 vss Q2 nCLK CLK DFlipFlop
.ends


* expanding   symbol:  mux2to4.sym # of pins=10
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/mux2to4.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/mux2to4.sch
.subckt mux2to4  vdd vss in_a in_b out_b_0 out_a_0 selec_0 out_b_1 out_a_1 selec_0_neg
*.iopin in_a
*.iopin in_b
*.ipin selec_0_neg
*.ipin selec_0
*.iopin out_b_0
*.iopin out_b_1
*.iopin out_a_0
*.iopin out_a_1
*.iopin vdd
*.iopin vss
x4 selec_0 out_a_1 in_a selec_0_neg vss vdd trans_gate_mux2to8
x5 selec_0_neg out_a_0 in_a selec_0 vss vdd trans_gate_mux2to8
x8 selec_0 out_b_1 in_b selec_0_neg vss vdd trans_gate_mux2to8
x9 selec_0_neg out_b_0 in_b selec_0 vss vdd trans_gate_mux2to8
.ends


* expanding   symbol:  mux2to1.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/mux2to1.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/mux2to1.sch
.subckt mux2to1  vdd vss in_a out_a_0 selec_0 out_a_1 selec_0_neg
*.iopin in_a
*.ipin selec_0_neg
*.ipin selec_0
*.iopin out_a_0
*.iopin out_a_1
*.iopin vdd
*.iopin vss
x4 selec_0 out_a_1 in_a selec_0_neg vss vdd trans_gate_mux2to8
x5 selec_0_neg out_a_0 in_a selec_0 vss vdd trans_gate_mux2to8
.ends


* expanding   symbol:  nor.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/nor.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/nor.sch
.subckt nor  vdd A B out vss
*.ipin A
*.ipin B
*.iopin vdd
*.opin out
*.iopin vss
XM1 out A vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out B vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 out B net1 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net1 A vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 net2 B vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 out A net2 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  inverter_csvco.sym # of pins=6
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_csvco.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_csvco.sch
.subckt inverter_csvco  vdd out in vss vbulkp vbulkn
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
*.iopin vbulkn
*.iopin vbulkp
XM1 out in vss vbulkn sky130_fd_pr__nfet_01v8 L=0.2 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out in vdd vbulkp sky130_fd_pr__pfet_01v8 L=0.2 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  latch_diff.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/latch_diff.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/latch_diff.sch
.subckt latch_diff  vdd nQ Q D nD CLK vss
*.iopin vdd
*.iopin vss
*.ipin D
*.opin nQ
*.ipin CLK
*.ipin nD
*.opin Q
XM3 net1 CLK vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM4 nQ Q vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM5 Q nQ vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM1 nQ D net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 Q nD net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:  mux_2to1_logic.sym # of pins=6
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/mux_2to1_logic.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/mux_2to1_logic.sch
.subckt mux_2to1_logic  avdd1p8 sel avss1p8 DinB out DinA
*.ipin DinB
*.ipin DinA
*.iopin avdd1p8
*.iopin avss1p8
*.ipin sel
*.opin out
XM5 out sel_b DinB avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=2.22 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM6 DinB sel out avss1p8 sky130_fd_pr__nfet_01v8 L=0.15 W=1.11 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out sel DinA avdd1p8 sky130_fd_pr__pfet_01v8 L=0.15 W=2.22 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7 DinA sel_b out avss1p8 sky130_fd_pr__nfet_01v8 L=0.15 W=1.11 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
x1 avdd1p8 sel_b sel avss1p8 inverter_min
.ends


* expanding   symbol:  buffer_no_inv_x05.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/buffer_no_inv_x05.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/buffer_no_inv_x05.sch
.subckt buffer_no_inv_x05  avdd1p8 in avss1p8 out
*.ipin in
*.iopin avdd1p8
*.iopin avss1p8
*.opin out
x1 avdd1p8 net1 in avss1p8 inverter_min
x2 avdd1p8 out net1 avss1p8 inverter_min
.ends


* expanding   symbol:  trans_gate_mux2to8.sym # of pins=6
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/trans_gate_mux2to8.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/trans_gate_mux2to8.sch
.subckt trans_gate_mux2to8  en_pos out in en_neg vss vdd
*.iopin en_neg
*.ipin in
*.opin out
*.iopin en_pos
*.iopin vdd
*.iopin vss
XM2 out en_neg in vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM1 out en_pos in vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
.ends


* expanding   symbol:  inverter_min.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_min.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_min.sch
.subckt inverter_min  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

** flattened .save nodes
.end
