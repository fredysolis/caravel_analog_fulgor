magic
tech sky130A
magscale 1 2
timestamp 1623892191
<< pwell >>
rect -2133 -2890 2133 2890
<< psubdiff >>
rect -2097 2820 -2001 2854
rect 2001 2820 2097 2854
rect -2097 2758 -2063 2820
rect 2063 2758 2097 2820
rect -2097 -2820 -2063 -2758
rect 2063 -2820 2097 -2758
rect -2097 -2854 -2001 -2820
rect 2001 -2854 2097 -2820
<< psubdiffcont >>
rect -2001 2820 2001 2854
rect -2097 -2758 -2063 2758
rect 2063 -2758 2097 2758
rect -2001 -2854 2001 -2820
<< xpolycontact >>
rect -1967 2292 -821 2724
rect -1967 -2724 -821 -2292
rect -573 2292 573 2724
rect -573 -2724 573 -2292
rect 821 2292 1967 2724
rect 821 -2724 1967 -2292
<< ppolyres >>
rect -1967 -2292 -821 2292
rect -573 -2292 573 2292
rect 821 -2292 1967 2292
<< locali >>
rect -2097 2820 -2001 2854
rect 2001 2820 2097 2854
rect -2097 2758 -2063 2820
rect 2063 2758 2097 2820
rect -2097 -2820 -2063 -2758
rect 2063 -2820 2097 -2758
rect -2097 -2854 -2001 -2820
rect 2001 -2854 2097 -2820
<< viali >>
rect -1951 2309 -837 2706
rect -557 2309 557 2706
rect 837 2309 1951 2706
rect -1951 -2706 -837 -2309
rect -557 -2706 557 -2309
rect 837 -2706 1951 -2309
<< metal1 >>
rect -1963 2706 -825 2712
rect -1963 2309 -1951 2706
rect -837 2309 -825 2706
rect -1963 2303 -825 2309
rect -569 2706 569 2712
rect -569 2309 -557 2706
rect 557 2309 569 2706
rect -569 2303 569 2309
rect 825 2706 1963 2712
rect 825 2309 837 2706
rect 1951 2309 1963 2706
rect 825 2303 1963 2309
rect -1963 -2309 -825 -2303
rect -1963 -2706 -1951 -2309
rect -837 -2706 -825 -2309
rect -1963 -2712 -825 -2706
rect -569 -2309 569 -2303
rect -569 -2706 -557 -2309
rect 557 -2706 569 -2309
rect -569 -2712 569 -2706
rect 825 -2309 1963 -2303
rect 825 -2706 837 -2309
rect 1951 -2706 1963 -2309
rect 825 -2712 1963 -2706
<< res5p73 >>
rect -1969 -2294 -819 2294
rect -575 -2294 575 2294
rect 819 -2294 1969 2294
<< properties >>
string gencell sky130_fd_pr__res_high_po_5p73
string FIXED_BBOX -2080 -2837 2080 2837
string parameters w 5.730 l 22.92 m 1 nx 3 wmin 5.730 lmin 0.50 rho 319.8 val 1.285k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 5.730 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
