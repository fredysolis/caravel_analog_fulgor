magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect -1127 -369 1127 369
<< pmos >>
rect -927 -150 -897 150
rect -831 -150 -801 150
rect -735 -150 -705 150
rect -639 -150 -609 150
rect -543 -150 -513 150
rect -447 -150 -417 150
rect -351 -150 -321 150
rect -255 -150 -225 150
rect -159 -150 -129 150
rect -63 -150 -33 150
rect 33 -150 63 150
rect 129 -150 159 150
rect 225 -150 255 150
rect 321 -150 351 150
rect 417 -150 447 150
rect 513 -150 543 150
rect 609 -150 639 150
rect 705 -150 735 150
rect 801 -150 831 150
rect 897 -150 927 150
<< pdiff >>
rect -989 138 -927 150
rect -989 -138 -977 138
rect -943 -138 -927 138
rect -989 -150 -927 -138
rect -897 138 -831 150
rect -897 -138 -881 138
rect -847 -138 -831 138
rect -897 -150 -831 -138
rect -801 138 -735 150
rect -801 -138 -785 138
rect -751 -138 -735 138
rect -801 -150 -735 -138
rect -705 138 -639 150
rect -705 -138 -689 138
rect -655 -138 -639 138
rect -705 -150 -639 -138
rect -609 138 -543 150
rect -609 -138 -593 138
rect -559 -138 -543 138
rect -609 -150 -543 -138
rect -513 138 -447 150
rect -513 -138 -497 138
rect -463 -138 -447 138
rect -513 -150 -447 -138
rect -417 138 -351 150
rect -417 -138 -401 138
rect -367 -138 -351 138
rect -417 -150 -351 -138
rect -321 138 -255 150
rect -321 -138 -305 138
rect -271 -138 -255 138
rect -321 -150 -255 -138
rect -225 138 -159 150
rect -225 -138 -209 138
rect -175 -138 -159 138
rect -225 -150 -159 -138
rect -129 138 -63 150
rect -129 -138 -113 138
rect -79 -138 -63 138
rect -129 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 129 150
rect 63 -138 79 138
rect 113 -138 129 138
rect 63 -150 129 -138
rect 159 138 225 150
rect 159 -138 175 138
rect 209 -138 225 138
rect 159 -150 225 -138
rect 255 138 321 150
rect 255 -138 271 138
rect 305 -138 321 138
rect 255 -150 321 -138
rect 351 138 417 150
rect 351 -138 367 138
rect 401 -138 417 138
rect 351 -150 417 -138
rect 447 138 513 150
rect 447 -138 463 138
rect 497 -138 513 138
rect 447 -150 513 -138
rect 543 138 609 150
rect 543 -138 559 138
rect 593 -138 609 138
rect 543 -150 609 -138
rect 639 138 705 150
rect 639 -138 655 138
rect 689 -138 705 138
rect 639 -150 705 -138
rect 735 138 801 150
rect 735 -138 751 138
rect 785 -138 801 138
rect 735 -150 801 -138
rect 831 138 897 150
rect 831 -138 847 138
rect 881 -138 897 138
rect 831 -150 897 -138
rect 927 138 989 150
rect 927 -138 943 138
rect 977 -138 989 138
rect 927 -150 989 -138
<< pdiffc >>
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
<< nsubdiff >>
rect -1057 299 -995 333
rect 995 299 1057 333
<< nsubdiffcont >>
rect -995 299 995 333
<< poly >>
rect -927 150 -897 176
rect -831 150 -801 176
rect -735 150 -705 176
rect -639 150 -609 176
rect -543 150 -513 176
rect -447 150 -417 176
rect -351 150 -321 176
rect -255 150 -225 176
rect -159 150 -129 176
rect -63 150 -33 176
rect 33 150 63 176
rect 129 150 159 176
rect 225 150 255 176
rect 321 150 351 176
rect 417 150 447 176
rect 513 150 543 176
rect 609 150 639 176
rect 705 150 735 176
rect 801 150 831 176
rect 897 150 927 176
rect -927 -181 -897 -150
rect -831 -181 -801 -150
rect -735 -181 -705 -150
rect -639 -181 -609 -150
rect -543 -181 -513 -150
rect -447 -181 -417 -150
rect -351 -181 -321 -150
rect -255 -181 -225 -150
rect -159 -181 -129 -150
rect -63 -181 -33 -150
rect -927 -247 -33 -181
rect 33 -181 63 -150
rect 129 -181 159 -150
rect 225 -181 255 -150
rect 321 -181 351 -150
rect 417 -181 447 -150
rect 513 -181 543 -150
rect 609 -181 639 -150
rect 705 -181 735 -150
rect 801 -181 831 -150
rect 897 -181 927 -150
rect 33 -247 927 -181
<< locali >>
rect -1057 299 -995 333
rect 995 299 1057 333
rect -977 138 -943 154
rect -977 -154 -943 -138
rect -881 138 -847 154
rect -881 -154 -847 -138
rect -785 138 -751 154
rect -785 -154 -751 -138
rect -689 138 -655 154
rect -689 -154 -655 -138
rect -593 138 -559 154
rect -593 -154 -559 -138
rect -497 138 -463 154
rect -497 -154 -463 -138
rect -401 138 -367 154
rect -401 -154 -367 -138
rect -305 138 -271 154
rect -305 -154 -271 -138
rect -209 138 -175 154
rect -209 -154 -175 -138
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect 175 138 209 154
rect 175 -154 209 -138
rect 271 138 305 154
rect 271 -154 305 -138
rect 367 138 401 154
rect 367 -154 401 -138
rect 463 138 497 154
rect 463 -154 497 -138
rect 559 138 593 154
rect 559 -154 593 -138
rect 655 138 689 154
rect 655 -154 689 -138
rect 751 138 785 154
rect 751 -154 785 -138
rect 847 138 881 154
rect 847 -154 881 -138
rect 943 138 977 154
rect 943 -154 977 -138
<< viali >>
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
<< metal1 >>
rect -983 138 -937 150
rect -983 -138 -977 138
rect -943 -138 -937 138
rect -983 -150 -937 -138
rect -887 138 -841 150
rect -887 -138 -881 138
rect -847 -138 -841 138
rect -887 -150 -841 -138
rect -791 138 -745 150
rect -791 -138 -785 138
rect -751 -138 -745 138
rect -791 -150 -745 -138
rect -695 138 -649 150
rect -695 -138 -689 138
rect -655 -138 -649 138
rect -695 -150 -649 -138
rect -599 138 -553 150
rect -599 -138 -593 138
rect -559 -138 -553 138
rect -599 -150 -553 -138
rect -503 138 -457 150
rect -503 -138 -497 138
rect -463 -138 -457 138
rect -503 -150 -457 -138
rect -407 138 -361 150
rect -407 -138 -401 138
rect -367 -138 -361 138
rect -407 -150 -361 -138
rect -311 138 -265 150
rect -311 -138 -305 138
rect -271 -138 -265 138
rect -311 -150 -265 -138
rect -215 138 -169 150
rect -215 -138 -209 138
rect -175 -138 -169 138
rect -215 -150 -169 -138
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -150 -73 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -150 119 -138
rect 169 138 215 150
rect 169 -138 175 138
rect 209 -138 215 138
rect 169 -150 215 -138
rect 265 138 311 150
rect 265 -138 271 138
rect 305 -138 311 138
rect 265 -150 311 -138
rect 361 138 407 150
rect 361 -138 367 138
rect 401 -138 407 138
rect 361 -150 407 -138
rect 457 138 503 150
rect 457 -138 463 138
rect 497 -138 503 138
rect 457 -150 503 -138
rect 553 138 599 150
rect 553 -138 559 138
rect 593 -138 599 138
rect 553 -150 599 -138
rect 649 138 695 150
rect 649 -138 655 138
rect 689 -138 695 138
rect 649 -150 695 -138
rect 745 138 791 150
rect 745 -138 751 138
rect 785 -138 791 138
rect 745 -150 791 -138
rect 841 138 887 150
rect 841 -138 847 138
rect 881 -138 887 138
rect 841 -150 887 -138
rect 937 138 983 150
rect 937 -138 943 138
rect 977 -138 983 138
rect 937 -150 983 -138
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1074 -316 1074 316
string parameters w 1.5 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
