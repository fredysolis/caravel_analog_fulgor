magic
tech sky130A
magscale 1 2
timestamp 1623893910
<< pwell >>
rect -16462 -24206 34360 5780
<< psubdiff >>
rect -16450 4360 -14850 4384
rect 32749 4360 34349 4384
rect 151 -145 175 -79
rect 4035 -145 4059 -79
rect -16450 -21664 -14850 -21640
rect -16450 -22594 -14851 -21664
rect 32749 -22593 34349 -21640
rect 32749 -22594 34348 -22593
rect -16450 -24194 -11039 -22594
rect 28961 -24194 34348 -22594
<< psubdiffcont >>
rect -16450 -21640 -14850 4360
rect 175 -145 4035 -79
rect 32749 -21640 34349 4360
rect -11039 -24194 28961 -22594
<< locali >>
rect -16450 4360 -14850 4376
rect 32749 4360 34349 4376
rect -14851 -21656 -14850 -21640
rect 34348 -21656 34349 -21640
<< viali >>
rect -16450 -21640 -14850 4360
rect 36 36 4230 70
rect 36 -79 4224 -49
rect 36 -145 175 -79
rect 175 -145 4035 -79
rect 4035 -145 4224 -79
rect 36 -168 4224 -145
rect -16450 -22594 -14851 -21640
rect 32749 -21640 34349 4360
rect 32749 -22594 34348 -21640
rect -16450 -24194 -11039 -22594
rect -11039 -24194 28961 -22594
rect 28961 -24194 34348 -22594
<< metal1 >>
rect -370 5080 -360 5680
rect 640 5614 650 5680
rect 2456 5614 2466 5680
rect 640 5182 1312 5614
rect 1560 5182 2466 5614
rect 640 5080 650 5182
rect 2456 5080 2466 5182
rect 3866 5614 3876 5680
rect 3866 5182 4100 5614
rect 3866 5080 3876 5182
rect -16456 4360 -14844 4372
rect -16456 -21634 -16450 4360
rect -16462 -24194 -16450 -21634
rect -14850 -21634 -14844 4360
rect 32743 4360 34355 4372
rect 166 166 3245 598
rect -10 70 4297 90
rect -10 36 36 70
rect 4230 36 4297 70
rect -10 -49 4297 36
rect -10 -168 36 -49
rect 4224 -168 4297 -49
rect -10 -185 4297 -168
rect 1312 -1221 2954 -185
rect 1312 -1273 2955 -1221
rect 1313 -2326 2955 -1273
rect -14850 -21640 -14839 -21634
rect -14851 -22588 -14839 -21640
rect 1313 -22588 2954 -2326
rect 32743 -22588 32749 4360
rect 34349 -21640 34355 4360
rect -14851 -22594 32749 -22588
rect 34348 -21652 34355 -21640
rect 34348 -22588 34354 -21652
rect 34348 -24194 34360 -22588
rect -16462 -24200 34360 -24194
rect 32743 -24206 34354 -24200
<< via1 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -10029 -23953 -4329 -22753
rect 9433 -24034 31413 -22834
<< metal2 >>
rect -360 5680 640 5690
rect -360 5070 640 5080
rect 2466 5680 3866 5690
rect 2466 5070 3866 5080
rect -10029 -22753 -4329 -22743
rect -10029 -23963 -4329 -23953
rect 9433 -22834 31413 -22824
rect 9433 -24044 31413 -24034
<< via2 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -10029 -23953 -4329 -22753
rect 9433 -24034 31413 -22834
<< metal3 >>
rect -370 5680 650 5685
rect -370 5080 -360 5680
rect 640 5080 650 5680
rect -370 5075 650 5080
rect 2456 5680 3876 5685
rect 2456 5080 2466 5680
rect 3866 5080 3876 5680
rect 2456 5075 3876 5080
rect -13523 -8002 -586 4898
rect -10029 -22748 -8629 -8002
rect -5695 -22748 -4295 -8002
rect 4852 -21602 31427 4898
rect -10039 -22753 -4295 -22748
rect -10039 -23953 -10029 -22753
rect -4329 -23136 -4295 -22753
rect 9433 -22829 10833 -21602
rect 14842 -22829 16242 -21602
rect 20055 -22829 21455 -21602
rect 25394 -22829 26794 -21602
rect 30027 -22829 31427 -21602
rect 9423 -22834 31427 -22829
rect -4329 -23953 -4319 -23136
rect -10039 -23958 -4319 -23953
rect 9423 -24034 9433 -22834
rect 31413 -23602 31427 -22834
rect 31413 -24034 31423 -23602
rect 9423 -24039 31423 -24034
rect 25394 -24061 26794 -24039
<< via3 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
<< metal4 >>
rect -12154 5680 740 5780
rect -12154 5080 -360 5680
rect 640 5080 740 5680
rect -12154 4980 740 5080
rect 2066 5680 29520 5780
rect 2066 5080 2466 5680
rect 3866 5080 29520 5680
rect 2066 4980 29520 5080
rect -12154 -6696 -10754 4980
rect -7779 -6696 -6379 4980
rect -3405 -6534 -2005 4980
rect 6722 -19031 8122 4980
rect 12166 -19023 13566 4980
rect 17484 -19174 18884 4980
rect 22862 -19265 24262 4980
rect 28119 -19235 29519 4980
use sky130_fd_pr__cap_mim_m3_1_W3JTNJ  sky130_fd_pr__cap_mim_m3_1_W3JTNJ_0
timestamp 1623892191
transform 1 0 -7054 0 1 -1552
box -6469 -6450 6468 6450
use sky130_fd_pr__cap_mim_m3_1_MA89VW  sky130_fd_pr__cap_mim_m3_1_MA89VW_0
timestamp 1623892191
transform 1 0 18140 0 1 -8352
box -13288 -13250 13287 13250
use sky130_fd_pr__res_high_po_5p73_GW5RGE  sky130_fd_pr__res_high_po_5p73_GW5RGE_0
timestamp 1623892191
transform 1 0 2133 0 1 2890
box -2133 -2890 2133 2890
<< labels >>
rlabel metal4 3866 4980 29520 5780 1 vc_pex
rlabel metal4 -12154 4980 -360 5780 1 in
rlabel metal1 1313 -22594 2954 -168 1 vss
<< end >>
