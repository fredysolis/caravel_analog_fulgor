magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect -455 -344 455 344
<< pmos >>
rect -255 -125 -225 125
rect -159 -125 -129 125
rect -63 -125 -33 125
rect 33 -125 63 125
rect 129 -125 159 125
rect 225 -125 255 125
<< pdiff >>
rect -317 113 -255 125
rect -317 -113 -305 113
rect -271 -113 -255 113
rect -317 -125 -255 -113
rect -225 113 -159 125
rect -225 -113 -209 113
rect -175 -113 -159 113
rect -225 -125 -159 -113
rect -129 113 -63 125
rect -129 -113 -113 113
rect -79 -113 -63 113
rect -129 -125 -63 -113
rect -33 113 33 125
rect -33 -113 -17 113
rect 17 -113 33 113
rect -33 -125 33 -113
rect 63 113 129 125
rect 63 -113 79 113
rect 113 -113 129 113
rect 63 -125 129 -113
rect 159 113 225 125
rect 159 -113 175 113
rect 209 -113 225 113
rect 159 -125 225 -113
rect 255 113 317 125
rect 255 -113 271 113
rect 305 -113 317 113
rect 255 -125 317 -113
<< pdiffc >>
rect -305 -113 -271 113
rect -209 -113 -175 113
rect -113 -113 -79 113
rect -17 -113 17 113
rect 79 -113 113 113
rect 175 -113 209 113
rect 271 -113 305 113
<< nsubdiff >>
rect -419 274 -323 308
rect 323 274 419 308
rect -419 212 -385 274
rect 385 212 419 274
rect -419 -274 -385 -212
rect 385 -274 419 -212
<< nsubdiffcont >>
rect -323 274 323 308
rect -419 -212 -385 212
rect 385 -212 419 212
<< poly >>
rect -255 125 -225 151
rect -159 125 -129 151
rect -63 125 -33 151
rect 33 125 63 151
rect 129 125 159 151
rect 225 125 255 151
rect -255 -154 -225 -125
rect -159 -154 -129 -125
rect -63 -154 -33 -125
rect 33 -154 63 -125
rect 129 -154 159 -125
rect 225 -154 255 -125
<< locali >>
rect -419 274 -323 308
rect 323 274 419 308
rect -419 212 -385 274
rect 385 212 419 274
rect -305 113 -271 129
rect -305 -129 -271 -113
rect -209 113 -175 129
rect -209 -129 -175 -113
rect -113 113 -79 129
rect -113 -129 -79 -113
rect -17 113 17 129
rect -17 -129 17 -113
rect 79 113 113 129
rect 79 -129 113 -113
rect 175 113 209 129
rect 175 -129 209 -113
rect 271 113 305 129
rect 271 -129 305 -113
rect -419 -274 -385 -212
rect 385 -274 419 -212
<< viali >>
rect -305 -113 -271 113
rect -209 -113 -175 113
rect -113 -113 -79 113
rect -17 -113 17 113
rect 79 -113 113 113
rect 175 -113 209 113
rect 271 -113 305 113
<< metal1 >>
rect -311 113 -265 125
rect -311 -113 -305 113
rect -271 -113 -265 113
rect -311 -125 -265 -113
rect -215 113 -169 125
rect -215 -113 -209 113
rect -175 -113 -169 113
rect -215 -125 -169 -113
rect -119 113 -73 125
rect -119 -113 -113 113
rect -79 -113 -73 113
rect -119 -125 -73 -113
rect -23 113 23 125
rect -23 -113 -17 113
rect 17 -113 23 113
rect -23 -125 23 -113
rect 73 113 119 125
rect 73 -113 79 113
rect 113 -113 119 113
rect 73 -125 119 -113
rect 169 113 215 125
rect 169 -113 175 113
rect 209 -113 215 113
rect 169 -125 215 -113
rect 265 113 311 125
rect 265 -113 271 113
rect 305 -113 311 113
rect 265 -125 311 -113
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -402 -291 402 291
string parameters w 1.25 l 0.15 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
