magic
tech sky130A
magscale 1 2
timestamp 1624395098
<< nwell >>
rect 3636 6239 4733 7015
rect 7538 6935 8332 7015
rect 7509 6239 7622 6935
rect 3666 4188 4554 4723
rect 3666 4000 4596 4188
rect 3666 3954 5436 4000
rect 3666 3947 7206 3954
rect 7538 3947 8332 4723
rect 3666 3890 8332 3947
rect 3666 3223 3976 3890
rect 3665 3206 3976 3223
rect 4556 3208 8332 3890
rect 4553 3206 8332 3208
rect 3665 3171 3959 3206
rect 4553 3171 4718 3206
rect 5436 3171 8332 3206
rect 3638 966 4062 1655
rect 6650 966 8332 1655
rect 3638 877 8332 966
rect 4054 871 8332 877
rect 6650 103 8332 871
rect 6650 -2189 8332 -1413
<< pwell >>
rect 3530 6050 4560 6239
rect 3530 5585 4978 6050
rect 3666 4723 4978 5585
rect 7389 5565 8332 6239
rect 7538 4723 8332 5565
rect 6650 2748 8332 3171
rect 3666 1655 8332 2748
rect 6650 -1413 8332 103
<< metal1 >>
rect 682 6891 736 6945
rect 3666 6851 4554 6985
rect 7538 6851 8332 6985
rect 3732 6209 3742 6289
rect 3985 6209 3995 6289
rect 4283 6195 4293 6273
rect 4460 6195 4470 6273
rect 7604 6199 7614 6284
rect 7857 6199 7867 6284
rect 8155 6195 8165 6273
rect 8332 6195 8342 6273
rect 2657 6067 2667 6121
rect 2926 6067 2936 6121
rect 6529 6074 6539 6130
rect 6798 6074 6808 6130
rect 3603 5645 4554 5813
rect 3666 5317 4554 5645
rect 7469 5317 8332 5813
rect 2651 4842 2661 4895
rect 2925 4842 2935 4895
rect 6523 4838 6533 4891
rect 6797 4838 6807 4891
rect 682 3977 754 3983
rect 3666 3981 4781 4111
rect 7195 3981 8332 4111
rect 3666 3977 8332 3981
rect 682 3917 8332 3977
rect 682 3911 754 3917
rect 3661 3783 8332 3917
rect 4556 3772 6572 3783
rect 4556 3737 4734 3772
rect 5432 3737 6572 3772
rect 7195 3701 8332 3783
rect 4025 3126 4035 3217
rect 4141 3126 4151 3217
rect 4236 3182 4246 3262
rect 4348 3182 4358 3262
rect 4436 3131 4798 3211
rect 5358 3127 5419 3205
rect 5556 3127 5927 3205
rect 5994 3193 6004 3262
rect 6126 3193 6136 3262
rect 6217 3131 6568 3211
rect 7130 3142 7183 3188
rect 2657 2999 2667 3051
rect 2926 2999 2936 3051
rect 4718 2623 5436 2690
rect 4718 2610 6488 2623
rect 6650 2610 8332 2743
rect 4718 2509 8332 2610
rect 3666 2249 8332 2509
rect 4062 2212 8332 2249
rect 6650 2083 8332 2212
rect 2656 1775 2666 1827
rect 2925 1775 2935 1827
rect 4780 1695 5017 1699
rect 4103 1615 4113 1695
rect 4230 1615 4240 1695
rect 4688 1615 4801 1637
rect 6509 1621 6519 1699
rect 6641 1621 6651 1699
rect 682 992 842 1003
rect 3666 992 4073 1043
rect 6650 992 8332 1126
rect 682 847 8332 992
rect 682 843 842 847
rect 6650 715 8332 847
rect 2656 -69 2666 -17
rect 2925 -69 2935 -17
rect 5641 -69 5651 -17
rect 5910 -69 5920 -17
rect 6650 -819 8332 -491
rect 2657 -1293 2667 -1241
rect 2926 -1293 2936 -1241
rect 5640 -1293 5650 -1241
rect 5909 -1293 5919 -1241
rect 682 -2119 747 -2065
rect 6650 -2159 8332 -2025
<< via1 >>
rect 3742 6209 3985 6289
rect 4293 6195 4460 6273
rect 7614 6199 7857 6284
rect 8165 6195 8332 6273
rect 2667 6067 2926 6121
rect 6539 6074 6798 6130
rect 2661 4842 2925 4895
rect 6533 4838 6797 4891
rect 4035 3126 4141 3217
rect 4246 3182 4348 3262
rect 5419 3127 5556 3205
rect 6004 3193 6126 3262
rect 2667 2999 2926 3051
rect 2666 1775 2925 1827
rect 4113 1615 4230 1695
rect 6519 1621 6641 1699
rect 2666 -69 2925 -17
rect 5651 -69 5910 -17
rect 2667 -1293 2926 -1241
rect 5650 -1293 5909 -1241
<< metal2 >>
rect 4814 6749 8283 6821
rect 924 6587 4397 6659
rect 924 6247 996 6587
rect 3742 6292 3985 6299
rect 3405 6289 3985 6292
rect 3405 6233 3742 6289
rect 4325 6283 4397 6587
rect 3742 6199 3985 6209
rect 4293 6273 4460 6283
rect 2667 6131 2926 6141
rect 2667 6057 2926 6067
rect 3866 6064 3925 6199
rect 4814 6228 4886 6749
rect 5429 6568 6704 6627
rect 4293 6185 4460 6195
rect 5429 6064 5488 6568
rect 6645 6140 6704 6568
rect 7614 6292 7857 6294
rect 7282 6284 7857 6292
rect 7282 6233 7614 6284
rect 8211 6283 8283 6749
rect 7614 6189 7857 6199
rect 8165 6273 8332 6283
rect 8165 6185 8332 6195
rect 6539 6130 6798 6140
rect 6539 6064 6798 6074
rect 3866 6005 5488 6064
rect 2661 4895 2925 4905
rect 2661 4822 2925 4832
rect 6533 4891 6797 4901
rect 6533 4812 6797 4822
rect 930 4250 1002 4726
rect 514 4178 1002 4250
rect 516 150 585 4178
rect 7309 3757 7381 4512
rect 1497 3685 7381 3757
rect 1497 3474 1569 3685
rect 926 3402 1569 3474
rect 926 3178 998 3402
rect 6004 3272 6126 3282
rect 4246 3262 4348 3272
rect 4035 3224 4141 3227
rect 3402 3217 4145 3224
rect 3402 3165 4035 3217
rect 4141 3165 4145 3217
rect 4246 3172 4348 3182
rect 5419 3205 5556 3215
rect 4035 3116 4141 3126
rect 2667 3060 2926 3070
rect 2667 2989 2926 2999
rect 4260 2417 4319 3172
rect 3713 2358 4319 2417
rect 6004 3173 6126 3183
rect 5419 3117 5556 3127
rect 2666 1827 2925 1837
rect 2666 1755 2925 1765
rect 3713 350 3772 2358
rect 5419 2265 5477 3117
rect 3473 291 3772 350
rect 3916 2207 5477 2265
rect 3916 341 3974 2207
rect 4113 1695 4230 1705
rect 4113 1605 4230 1615
rect 6519 1699 6641 1709
rect 6519 1611 6641 1621
rect 4115 1016 4173 1605
rect 4115 958 6488 1016
rect 516 81 1027 150
rect 3916 118 3975 341
rect 6430 138 6488 958
rect 2666 -7 2925 3
rect 2666 -79 2925 -69
rect 5651 -7 5910 3
rect 5651 -79 5910 -69
rect 2667 -1241 2926 -1231
rect 2667 -1313 2926 -1303
rect 5650 -1241 5909 -1231
rect 5650 -1313 5909 -1303
<< via2 >>
rect 2667 6121 2926 6131
rect 2667 6067 2926 6121
rect 4293 6195 4460 6273
rect 8165 6195 8332 6273
rect 2661 4842 2925 4895
rect 2661 4832 2925 4842
rect 6533 4838 6797 4891
rect 6533 4822 6797 4838
rect 6004 3262 6126 3272
rect 2667 3051 2926 3060
rect 2667 2999 2926 3051
rect 6004 3193 6126 3262
rect 6004 3183 6126 3193
rect 2666 1775 2925 1827
rect 2666 1765 2925 1775
rect 2666 -17 2925 -7
rect 2666 -69 2925 -17
rect 5651 -17 5910 -7
rect 5651 -69 5910 -17
rect 2667 -1293 2926 -1241
rect 2667 -1303 2926 -1293
rect 5650 -1293 5909 -1241
rect 5650 -1303 5909 -1293
<< metal3 >>
rect 4283 6273 4470 6278
rect 4283 6195 4293 6273
rect 4460 6195 4470 6273
rect 4283 6190 4470 6195
rect 8155 6273 8342 6278
rect 8155 6195 8165 6273
rect 8332 6195 8342 6273
rect 8155 6190 8342 6195
rect 2657 6067 2667 6141
rect 2926 6067 2936 6141
rect 2657 6062 2936 6067
rect 2651 4895 2935 4900
rect 118 4821 128 4895
rect 228 4821 238 4895
rect 2651 4822 2661 4895
rect 2925 4822 2935 4895
rect 127 1828 228 4821
rect 4334 3898 4408 6190
rect 6523 4891 6807 4896
rect 6523 4822 6533 4891
rect 6797 4822 6807 4891
rect 6523 4817 6807 4822
rect 6683 3898 6757 4817
rect 4334 3824 6757 3898
rect 5994 3272 6136 3277
rect 5994 3183 6004 3272
rect 6126 3183 6136 3272
rect 5994 3178 6136 3183
rect 2657 2999 2667 3070
rect 2926 2999 2936 3070
rect 2657 2994 2936 2999
rect 118 1754 128 1828
rect 228 1754 238 1828
rect 2656 1827 2935 1832
rect 2656 1755 2666 1827
rect 2925 1755 2935 1827
rect 127 4 228 1754
rect 2684 1261 2758 1755
rect 6028 1261 6102 3178
rect 2684 1187 6102 1261
rect 117 -70 127 4
rect 228 -70 238 4
rect 2656 -69 2666 3
rect 2925 -69 2935 3
rect 2656 -74 2935 -69
rect 5641 -69 5651 3
rect 5910 -69 5920 3
rect 5641 -74 5920 -69
rect 2657 -1241 2936 -1236
rect 2657 -1313 2667 -1241
rect 2926 -1313 2936 -1241
rect 5640 -1241 5919 -1236
rect 5640 -1313 5650 -1241
rect 5909 -1313 5919 -1241
<< via3 >>
rect 2667 6131 2926 6141
rect 2667 6067 2926 6131
rect 128 4821 228 4895
rect 2661 4832 2925 4895
rect 2661 4822 2925 4832
rect 2667 3060 2926 3070
rect 2667 2999 2926 3060
rect 128 1754 228 1828
rect 2666 1765 2925 1827
rect 2666 1755 2925 1765
rect 127 -70 228 4
rect 2666 -7 2925 3
rect 2666 -69 2925 -7
rect 5651 -7 5910 3
rect 5651 -69 5910 -7
rect 2667 -1303 2926 -1241
rect 2667 -1313 2926 -1303
rect 5650 -1303 5909 -1241
rect 5650 -1313 5909 -1303
<< metal4 >>
rect 2666 6141 2927 6142
rect 2666 6140 2667 6141
rect -92 6067 2667 6140
rect 2926 6067 2927 6141
rect -92 6066 2927 6067
rect -92 3072 -18 6066
rect 127 4895 229 4896
rect 2660 4895 2926 4896
rect 127 4821 128 4895
rect 228 4822 2661 4895
rect 2925 4822 2926 4895
rect 228 4821 2926 4822
rect 127 4820 229 4821
rect -92 3071 2772 3072
rect -92 3070 2927 3071
rect -92 2999 2667 3070
rect 2926 2999 2927 3070
rect -92 2998 2927 2999
rect -92 -1240 -18 2998
rect 127 1828 229 1829
rect 127 1754 128 1828
rect 228 1827 2926 1828
rect 228 1755 2666 1827
rect 2925 1755 2926 1827
rect 228 1754 2926 1755
rect 127 1753 229 1754
rect 126 4 229 5
rect 126 -70 127 4
rect 228 3 5911 4
rect 228 -69 2666 3
rect 2925 -69 5651 3
rect 5910 -69 5911 3
rect 228 -70 5911 -69
rect 126 -71 229 -70
rect -92 -1241 5910 -1240
rect -92 -1313 2667 -1241
rect 2926 -1313 5650 -1241
rect 5909 -1313 5910 -1241
rect -92 -1314 5910 -1313
use DFlipFlop  DFlipFlop_2
timestamp 1624049879
transform 1 0 1926 0 1 879
box -1244 0 1740 3068
use DFlipFlop  DFlipFlop_3
timestamp 1624049879
transform 1 0 1926 0 -1 879
box -1244 0 1740 3068
use DFlipFlop  DFlipFlop_4
timestamp 1624049879
transform 1 0 4910 0 -1 879
box -1244 0 1740 3068
use nand_logic  nand_logic_0
timestamp 1623952422
transform 1 0 3885 0 1 3205
box -219 -731 833 707
use DFlipFlop  DFlipFlop_0
timestamp 1624049879
transform 1 0 1926 0 1 3947
box -1244 0 1740 3068
use inverter_min_x16  inverter_min_x16_0
timestamp 1624046389
transform 1 0 4833 0 -1 1602
box -53 -616 1817 643
use nand_logic  nand_logic_1
timestamp 1623952422
transform 1 0 5655 0 1 3205
box -219 -731 833 707
use inverter_min_x4  inverter_min_x4_1
timestamp 1624049879
transform 1 0 4771 0 1 3224
box -53 -616 665 643
use inverter_min_x4  inverter_min_x4_3
timestamp 1624049879
transform 1 0 6541 0 1 3224
box -53 -616 665 643
use inverter_min_x4  inverter_min_x4_4
timestamp 1624049879
transform 1 0 4115 0 -1 1602
box -53 -616 665 643
use DFlipFlop  DFlipFlop_1
timestamp 1624049879
transform 1 0 5798 0 1 3947
box -1244 0 1740 3068
use inverter_min_x4  inverter_min_x4_0
timestamp 1624049879
transform 1 0 3795 0 1 6292
box -53 -616 665 643
use inverter_min_x4  inverter_min_x4_2
timestamp 1624049879
transform 1 0 7667 0 1 6292
box -53 -616 665 643
<< labels >>
rlabel metal1 7614 5716 8332 5771 1 vss
rlabel metal1 7469 5317 7538 5645 5 vss
rlabel via1 6551 1642 6601 1680 1 clk_amp
rlabel metal4 -64 -38 -36 -5 1 clkn
rlabel metal1 702 6909 718 6931 1 avdd1p8
rlabel metal1 7130 3142 7183 3188 1 rst
rlabel metal3 159 4649 206 4710 1 clkp
rlabel metal1 7948 5421 8048 5515 1 avss1p8
rlabel metal1 7873 2391 7973 2485 1 avss1p8
rlabel metal1 7805 -720 7905 -626 1 avss1p8
<< end >>
