**.subckt top_pll_v1_pex_no_integration vdd vss in_ref pfd_QA pfd_QB Up nUp Down nDown pfd_reset
*+ cp_nswitch cp_pswitch cp_biasp iref_cp lf_vc D0_vco vco_vctrl vco_out out_first_buffer out_to_pad out_to_div
*+ out_by_2 n_out_by_2 out_div_2 n_out_div_2 out_buffer_div_2 n_out_buffer_div_2 div_5_Q1 div_5_Q1_shift
*+ div_5_nQ0 div_5_Q0 div_5_nQ2 out_div_by_5 out_to_buffer D0_cap
*.iopin vdd
*.iopin vss
*.ipin in_ref
*.iopin pfd_QA
*.iopin pfd_QB
*.iopin Up
*.iopin nUp
*.iopin Down
*.iopin nDown
*.iopin pfd_reset
*.iopin cp_nswitch
*.iopin cp_pswitch
*.iopin cp_biasp
*.ipin iref_cp
*.iopin lf_vc
*.iopin D0_vco
*.iopin vco_vctrl
*.iopin vco_out
*.iopin out_first_buffer
*.opin out_to_pad
*.iopin out_to_div
*.iopin out_by_2
*.iopin n_out_by_2
*.iopin out_div_2
*.iopin n_out_div_2
*.iopin out_buffer_div_2
*.iopin n_out_buffer_div_2
*.iopin div_5_Q1
*.iopin div_5_Q1_shift
*.iopin div_5_nQ0
*.iopin div_5_Q0
*.iopin div_5_nQ2
*.iopin out_div_by_5
*.iopin out_to_buffer
*.iopin D0_cap
x1 vss vdd pfd_QA in_ref out_div_by_5 pfd_QB pfd_reset PFD_pex_c
x2 vdd Up nUp vco_vctrl Down nDown vss iref_cp cp_nswitch cp_pswitch cp_biasp charge_pump_pex_c
x3 vdd vco_out vco_vctrl vss D0_vco csvco_pex_c
x5 vdd out_div_by_5 out_by_2 vss n_out_by_2 div_5_nQ2 div_5_Q1 div_5_nQ0 div_5_Q0 div_5_Q1_shift
+ div_by_5_pex_c
x7 Up vdd pfd_QA nUp Down pfd_QB vss nDown pfd_cp_interface_pex_c
x8 vdd vco_out out_to_buffer out_to_div vss out_first_buffer ring_osc_buffer_pex_c
x4 n_out_by_2 vss out_to_div vdd out_by_2 out_div_2 n_out_div_2 out_buffer_div_2 n_out_buffer_div_2
+ div_by_2_pex_c
x9 vdd out_to_pad out_to_buffer vss buffer_salida_pex_c
x6 vss vco_vctrl lf_vc D0_cap loop_filter_v2
**.ends

* expanding   symbol:  loop_filter_v2.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/loop_filter_v2.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/loop_filter_v2.sch
.subckt loop_filter_v2  vss in vc_pex D0_cap
*.iopin in
*.iopin vss
*.iopin vc_pex
*.iopin D0_cap
x1 in net1 vss res_loop_filter
x2 vc_pex net1 vss res_loop_filter
x3 vc_pex net1 vss res_loop_filter
x4 vc_pex vss cap1_loop_filter
x5 in vss cap2_loop_filter
XM1 in D0_cap net2 vss sky130_fd_pr__nfet_01v8 L=0.3 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x6 net2 vss cap3_loop_filter
.ends


* expanding   symbol:  res_loop_filter.sym # of pins=3
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/res_loop_filter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/res_loop_filter.sch
.subckt res_loop_filter  in out vss
*.iopin in
*.iopin vss
*.iopin out
XR3 out in vss sky130_fd_pr__res_high_po_5p73 L=22.92 mult=1 m=1
.ends


* expanding   symbol:  cap1_loop_filter.sym # of pins=2
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/cap1_loop_filter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/cap1_loop_filter.sch
.subckt cap1_loop_filter  in out
*.iopin in
*.iopin out
XC1 in out sky130_fd_pr__cap_mim_m3_1 W=25 L=25 MF=25 m=25
.ends


* expanding   symbol:  cap2_loop_filter.sym # of pins=2
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/cap2_loop_filter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/cap2_loop_filter.sch
.subckt cap2_loop_filter  in out
*.iopin in
*.iopin out
XC1 in out sky130_fd_pr__cap_mim_m3_1 W=20 L=20 MF=9 m=9
.ends


* expanding   symbol:  cap3_loop_filter.sym # of pins=2
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/cap3_loop_filter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/cap3_loop_filter.sch
.subckt cap3_loop_filter  in out
*.iopin in
*.iopin out
XC1 in out sky130_fd_pr__cap_mim_m3_1 W=20 L=20 MF=4 m=4
.ends

** flattened .save nodes
.end
