* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A


* Top level circuit user_analog_project_wrapper

.end

