magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect -2457 -634 2457 634
<< pmos >>
rect -2261 -486 -1861 414
rect -1803 -486 -1403 414
rect -1345 -486 -945 414
rect -887 -486 -487 414
rect -429 -486 -29 414
rect 29 -486 429 414
rect 487 -486 887 414
rect 945 -486 1345 414
rect 1403 -486 1803 414
rect 1861 -486 2261 414
<< pdiff >>
rect -2319 402 -2261 414
rect -2319 -474 -2307 402
rect -2273 -474 -2261 402
rect -2319 -486 -2261 -474
rect -1861 402 -1803 414
rect -1861 -474 -1849 402
rect -1815 -474 -1803 402
rect -1861 -486 -1803 -474
rect -1403 402 -1345 414
rect -1403 -474 -1391 402
rect -1357 -474 -1345 402
rect -1403 -486 -1345 -474
rect -945 402 -887 414
rect -945 -474 -933 402
rect -899 -474 -887 402
rect -945 -486 -887 -474
rect -487 402 -429 414
rect -487 -474 -475 402
rect -441 -474 -429 402
rect -487 -486 -429 -474
rect -29 402 29 414
rect -29 -474 -17 402
rect 17 -474 29 402
rect -29 -486 29 -474
rect 429 402 487 414
rect 429 -474 441 402
rect 475 -474 487 402
rect 429 -486 487 -474
rect 887 402 945 414
rect 887 -474 899 402
rect 933 -474 945 402
rect 887 -486 945 -474
rect 1345 402 1403 414
rect 1345 -474 1357 402
rect 1391 -474 1403 402
rect 1345 -486 1403 -474
rect 1803 402 1861 414
rect 1803 -474 1815 402
rect 1849 -474 1861 402
rect 1803 -486 1861 -474
rect 2261 402 2319 414
rect 2261 -474 2273 402
rect 2307 -474 2319 402
rect 2261 -486 2319 -474
<< pdiffc >>
rect -2307 -474 -2273 402
rect -1849 -474 -1815 402
rect -1391 -474 -1357 402
rect -933 -474 -899 402
rect -475 -474 -441 402
rect -17 -474 17 402
rect 441 -474 475 402
rect 899 -474 933 402
rect 1357 -474 1391 402
rect 1815 -474 1849 402
rect 2273 -474 2307 402
<< nsubdiff >>
rect -2387 -598 -2325 -564
rect 2325 -598 2387 -564
<< nsubdiffcont >>
rect -2325 -598 2325 -564
<< poly >>
rect -2261 455 2261 511
rect -2261 414 -1861 455
rect -1803 414 -1403 455
rect -1345 414 -945 455
rect -887 414 -487 455
rect -429 414 -29 455
rect 29 414 429 455
rect 487 414 887 455
rect 945 414 1345 455
rect 1403 414 1803 455
rect 1861 414 2261 455
rect -2261 -512 -1861 -486
rect -1803 -512 -1403 -486
rect -1345 -512 -945 -486
rect -887 -512 -487 -486
rect -429 -512 -29 -486
rect 29 -512 429 -486
rect 487 -512 887 -486
rect 945 -512 1345 -486
rect 1403 -512 1803 -486
rect 1861 -512 2261 -486
<< locali >>
rect -2307 402 -2273 418
rect -2307 -490 -2273 -474
rect -1849 402 -1815 418
rect -1849 -490 -1815 -474
rect -1391 402 -1357 418
rect -1391 -490 -1357 -474
rect -933 402 -899 418
rect -933 -490 -899 -474
rect -475 402 -441 418
rect -475 -490 -441 -474
rect -17 402 17 418
rect -17 -490 17 -474
rect 441 402 475 418
rect 441 -490 475 -474
rect 899 402 933 418
rect 899 -490 933 -474
rect 1357 402 1391 418
rect 1357 -490 1391 -474
rect 1815 402 1849 418
rect 1815 -490 1849 -474
rect 2273 402 2307 418
rect 2273 -490 2307 -474
rect -2387 -598 -2325 -564
rect 2325 -598 2387 -564
<< viali >>
rect -2307 -474 -2273 402
rect -1849 -474 -1815 402
rect -1391 -474 -1357 402
rect -933 -474 -899 402
rect -475 -474 -441 402
rect -17 -474 17 402
rect 441 -474 475 402
rect 899 -474 933 402
rect 1357 -474 1391 402
rect 1815 -474 1849 402
rect 2273 -474 2307 402
<< metal1 >>
rect -2313 402 -2267 414
rect -2313 -474 -2307 402
rect -2273 -474 -2267 402
rect -2313 -486 -2267 -474
rect -1855 402 -1809 414
rect -1855 -474 -1849 402
rect -1815 -474 -1809 402
rect -1855 -486 -1809 -474
rect -1397 402 -1351 414
rect -1397 -474 -1391 402
rect -1357 -474 -1351 402
rect -1397 -486 -1351 -474
rect -939 402 -893 414
rect -939 -474 -933 402
rect -899 -474 -893 402
rect -939 -486 -893 -474
rect -481 402 -435 414
rect -481 -474 -475 402
rect -441 -474 -435 402
rect -481 -486 -435 -474
rect -23 402 23 414
rect -23 -474 -17 402
rect 17 -474 23 402
rect -23 -486 23 -474
rect 435 402 481 414
rect 435 -474 441 402
rect 475 -474 481 402
rect 435 -486 481 -474
rect 893 402 939 414
rect 893 -474 899 402
rect 933 -474 939 402
rect 893 -486 939 -474
rect 1351 402 1397 414
rect 1351 -474 1357 402
rect 1391 -474 1397 402
rect 1351 -486 1397 -474
rect 1809 402 1855 414
rect 1809 -474 1815 402
rect 1849 -474 1855 402
rect 1809 -486 1855 -474
rect 2267 402 2313 414
rect 2267 -474 2273 402
rect 2307 -474 2313 402
rect 2267 -486 2313 -474
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -2404 -581 2404 581
string parameters w 4.5 l 2 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
