magic
tech sky130A
magscale 1 2
timestamp 1623774805
<< pwell >>
rect -1957 -254 1957 254
<< nmos >>
rect -1761 -44 -1461 106
rect -1403 -44 -1103 106
rect -1045 -44 -745 106
rect -687 -44 -387 106
rect -329 -44 -29 106
rect 29 -44 329 106
rect 387 -44 687 106
rect 745 -44 1045 106
rect 1103 -44 1403 106
rect 1461 -44 1761 106
<< ndiff >>
rect -1819 94 -1761 106
rect -1819 -32 -1807 94
rect -1773 -32 -1761 94
rect -1819 -44 -1761 -32
rect -1461 94 -1403 106
rect -1461 -32 -1449 94
rect -1415 -32 -1403 94
rect -1461 -44 -1403 -32
rect -1103 94 -1045 106
rect -1103 -32 -1091 94
rect -1057 -32 -1045 94
rect -1103 -44 -1045 -32
rect -745 94 -687 106
rect -745 -32 -733 94
rect -699 -32 -687 94
rect -745 -44 -687 -32
rect -387 94 -329 106
rect -387 -32 -375 94
rect -341 -32 -329 94
rect -387 -44 -329 -32
rect -29 94 29 106
rect -29 -32 -17 94
rect 17 -32 29 94
rect -29 -44 29 -32
rect 329 94 387 106
rect 329 -32 341 94
rect 375 -32 387 94
rect 329 -44 387 -32
rect 687 94 745 106
rect 687 -32 699 94
rect 733 -32 745 94
rect 687 -44 745 -32
rect 1045 94 1103 106
rect 1045 -32 1057 94
rect 1091 -32 1103 94
rect 1045 -44 1103 -32
rect 1403 94 1461 106
rect 1403 -32 1415 94
rect 1449 -32 1461 94
rect 1403 -44 1461 -32
rect 1761 94 1819 106
rect 1761 -32 1773 94
rect 1807 -32 1819 94
rect 1761 -44 1819 -32
<< ndiffc >>
rect -1807 -32 -1773 94
rect -1449 -32 -1415 94
rect -1091 -32 -1057 94
rect -733 -32 -699 94
rect -375 -32 -341 94
rect -17 -32 17 94
rect 341 -32 375 94
rect 699 -32 733 94
rect 1057 -32 1091 94
rect 1415 -32 1449 94
rect 1773 -32 1807 94
<< psubdiff >>
rect -1887 184 -1825 218
rect 1825 184 1887 218
<< psubdiffcont >>
rect -1825 184 1825 218
<< poly >>
rect -1761 106 -1461 132
rect -1403 106 -1103 132
rect -1045 106 -745 132
rect -687 106 -387 132
rect -329 106 -29 132
rect 29 106 329 132
rect 387 106 687 132
rect 745 106 1045 132
rect 1103 106 1403 132
rect 1461 106 1761 132
rect -1761 -66 -1461 -44
rect -1403 -66 -1103 -44
rect -1045 -66 -745 -44
rect -687 -66 -387 -44
rect -329 -66 -29 -44
rect 29 -66 329 -44
rect 387 -66 687 -44
rect 745 -66 1045 -44
rect 1103 -66 1403 -44
rect 1461 -66 1761 -44
rect -1761 -132 1761 -66
<< locali >>
rect -1887 184 -1825 218
rect 1825 184 1887 218
rect -1807 94 -1773 110
rect -1807 -48 -1773 -32
rect -1449 94 -1415 110
rect -1449 -48 -1415 -32
rect -1091 94 -1057 110
rect -1091 -48 -1057 -32
rect -733 94 -699 110
rect -733 -48 -699 -32
rect -375 94 -341 110
rect -375 -48 -341 -32
rect -17 94 17 110
rect -17 -48 17 -32
rect 341 94 375 110
rect 341 -48 375 -32
rect 699 94 733 110
rect 699 -48 733 -32
rect 1057 94 1091 110
rect 1057 -48 1091 -32
rect 1415 94 1449 110
rect 1415 -48 1449 -32
rect 1773 94 1807 110
rect 1773 -48 1807 -32
<< viali >>
rect -1807 -32 -1773 94
rect -1449 -32 -1415 94
rect -1091 -32 -1057 94
rect -733 -32 -699 94
rect -375 -32 -341 94
rect -17 -32 17 94
rect 341 -32 375 94
rect 699 -32 733 94
rect 1057 -32 1091 94
rect 1415 -32 1449 94
rect 1773 -32 1807 94
<< metal1 >>
rect -1813 94 -1767 106
rect -1813 -32 -1807 94
rect -1773 -32 -1767 94
rect -1813 -44 -1767 -32
rect -1455 94 -1409 106
rect -1455 -32 -1449 94
rect -1415 -32 -1409 94
rect -1455 -44 -1409 -32
rect -1097 94 -1051 106
rect -1097 -32 -1091 94
rect -1057 -32 -1051 94
rect -1097 -44 -1051 -32
rect -739 94 -693 106
rect -739 -32 -733 94
rect -699 -32 -693 94
rect -739 -44 -693 -32
rect -381 94 -335 106
rect -381 -32 -375 94
rect -341 -32 -335 94
rect -381 -44 -335 -32
rect -23 94 23 106
rect -23 -32 -17 94
rect 17 -32 23 94
rect -23 -44 23 -32
rect 335 94 381 106
rect 335 -32 341 94
rect 375 -32 381 94
rect 335 -44 381 -32
rect 693 94 739 106
rect 693 -32 699 94
rect 733 -32 739 94
rect 693 -44 739 -32
rect 1051 94 1097 106
rect 1051 -32 1057 94
rect 1091 -32 1097 94
rect 1051 -44 1097 -32
rect 1409 94 1455 106
rect 1409 -32 1415 94
rect 1449 -32 1455 94
rect 1409 -44 1455 -32
rect 1767 94 1813 106
rect 1767 -32 1773 94
rect 1807 -32 1813 94
rect 1767 -44 1813 -32
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1904 -201 1904 201
string parameters w 0.75 l 1.5 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
