magic
tech sky130A
magscale 1 2
timestamp 1623972527
<< nwell >>
rect -257 -702 257 701
<< pmos >>
rect -159 -600 -129 600
rect -63 -600 -33 600
rect 33 -600 63 600
rect 129 -600 159 600
<< pdiff >>
rect -221 588 -159 600
rect -221 -588 -209 588
rect -175 -588 -159 588
rect -221 -600 -159 -588
rect -129 588 -63 600
rect -129 -588 -113 588
rect -79 -588 -63 588
rect -129 -600 -63 -588
rect -33 588 33 600
rect -33 -588 -17 588
rect 17 -588 33 588
rect -33 -600 33 -588
rect 63 588 129 600
rect 63 -588 79 588
rect 113 -588 129 588
rect 63 -600 129 -588
rect 159 588 221 600
rect 159 -588 175 588
rect 209 -588 221 588
rect 159 -600 221 -588
<< pdiffc >>
rect -209 -588 -175 588
rect -113 -588 -79 588
rect -17 -588 17 588
rect 79 -588 113 588
rect 175 -588 209 588
<< poly >>
rect -257 624 257 695
rect -159 600 -129 624
rect -63 600 -33 624
rect 33 600 63 624
rect 129 600 159 624
rect -159 -621 -129 -600
rect -63 -621 -33 -600
rect 33 -621 63 -600
rect 129 -621 159 -600
rect -257 -777 257 -621
<< locali >>
rect -209 588 -175 604
rect -209 -604 -175 -588
rect -113 588 -79 604
rect -113 -604 -79 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 79 588 113 604
rect 79 -604 113 -588
rect 175 588 209 604
rect 175 -604 209 -588
<< viali >>
rect -209 -588 -175 588
rect -113 -588 -79 588
rect -17 -588 17 588
rect 79 -588 113 588
rect 175 -588 209 588
<< metal1 >>
rect -257 685 257 744
rect -215 588 -169 685
rect -215 -588 -209 588
rect -175 -588 -169 588
rect -215 -600 -169 -588
rect -119 588 -73 600
rect -119 -588 -113 588
rect -79 -588 -73 588
rect -119 -636 -73 -588
rect -23 588 23 685
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 73 588 119 600
rect 73 -588 79 588
rect 113 -588 119 588
rect 73 -636 119 -588
rect 169 588 215 685
rect 169 -588 175 588
rect 209 -588 215 588
rect 169 -600 215 -588
rect -257 -723 257 -636
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 6 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
