magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< metal3 >>
rect -42552 -37389 -15977 -16050
rect -42552 -37390 -35133 -37389
rect -42552 -37422 -40452 -37390
rect -39452 -37421 -35133 -37390
rect -34133 -37421 -29815 -37389
rect -28815 -37421 -24497 -37389
rect -23497 -37421 -19179 -37389
rect -18179 -37421 -15977 -37389
rect -39452 -37422 -15977 -37421
rect -42552 -40573 -15977 -37422
rect -42552 -42450 -16417 -40573
rect -40452 -42690 -39452 -42450
rect -35133 -42690 -34133 -42450
rect -29815 -42690 -28815 -42450
rect -24497 -42690 -23497 -42450
rect -19179 -42690 -18179 -42450
rect -17417 -42678 -16417 -42450
rect -40452 -43690 -18179 -42690
<< metal4 >>
rect -40452 -15842 -18179 -14842
rect -40452 -21110 -39452 -15842
rect -35133 -21111 -34133 -15842
rect -29815 -21111 -28815 -15842
rect -24497 -21111 -23497 -15842
rect -19179 -21111 -18179 -15842
use sky130_fd_pr__cap_mim_m3_1_MACBVW  sky130_fd_pr__cap_mim_m3_1_MACBVW_0
timestamp 1624049879
transform 1 0 -29264 0 1 -29250
box -13288 -13200 13287 13200
<< labels >>
rlabel metal4 -40452 -15842 -18179 -14842 1 in
rlabel metal3 -40452 -43690 -18179 -42690 1 out
<< end >>
