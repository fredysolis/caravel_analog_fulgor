magic
tech sky130A
magscale 1 2
timestamp 1624030292
<< nwell >>
rect -487 -419 487 419
<< pmoslvt >>
rect -291 -200 -221 200
rect -163 -200 -93 200
rect -35 -200 35 200
rect 93 -200 163 200
rect 221 -200 291 200
<< pdiff >>
rect -349 188 -291 200
rect -349 -188 -337 188
rect -303 -188 -291 188
rect -349 -200 -291 -188
rect -221 188 -163 200
rect -221 -188 -209 188
rect -175 -188 -163 188
rect -221 -200 -163 -188
rect -93 188 -35 200
rect -93 -188 -81 188
rect -47 -188 -35 188
rect -93 -200 -35 -188
rect 35 188 93 200
rect 35 -188 47 188
rect 81 -188 93 188
rect 35 -200 93 -188
rect 163 188 221 200
rect 163 -188 175 188
rect 209 -188 221 188
rect 163 -200 221 -188
rect 291 188 349 200
rect 291 -188 303 188
rect 337 -188 349 188
rect 291 -200 349 -188
<< pdiffc >>
rect -337 -188 -303 188
rect -209 -188 -175 188
rect -81 -188 -47 188
rect 47 -188 81 188
rect 175 -188 209 188
rect 303 -188 337 188
<< nsubdiff >>
rect -451 349 -355 383
rect 355 349 451 383
rect -451 287 -417 349
rect 417 287 451 349
rect -451 -349 -417 -287
rect 417 -349 451 -287
rect -451 -383 -355 -349
rect 355 -383 451 -349
<< nsubdiffcont >>
rect -355 349 355 383
rect -451 -287 -417 287
rect 417 -287 451 287
rect -355 -383 355 -349
<< poly >>
rect -291 281 291 297
rect -291 247 -275 281
rect -237 247 -147 281
rect -109 247 -19 281
rect 19 247 109 281
rect 147 247 237 281
rect 275 247 291 281
rect -291 233 291 247
rect -291 200 -221 233
rect -163 200 -93 233
rect -35 200 35 233
rect 93 200 163 233
rect 221 200 291 233
rect -291 -238 -221 -200
rect -163 -238 -93 -200
rect -35 -238 35 -200
rect 93 -238 163 -200
rect 221 -238 291 -200
<< polycont >>
rect -275 247 -237 281
rect -147 247 -109 281
rect -19 247 19 281
rect 109 247 147 281
rect 237 247 275 281
<< locali >>
rect -451 349 -355 383
rect 355 349 451 383
rect -451 287 -417 349
rect 417 287 451 349
rect -291 247 -275 281
rect 275 247 291 281
rect -337 188 -303 204
rect -337 -204 -303 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -81 188 -47 204
rect -81 -204 -47 -188
rect 47 188 81 204
rect 47 -204 81 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 303 188 337 204
rect 303 -204 337 -188
rect -451 -349 -417 -287
rect 417 -349 451 -287
rect -451 -383 -355 -349
rect 355 -383 451 -349
<< viali >>
rect -275 247 -237 281
rect -237 247 -147 281
rect -147 247 -109 281
rect -109 247 -19 281
rect -19 247 19 281
rect 19 247 109 281
rect 109 247 147 281
rect 147 247 237 281
rect 237 247 275 281
rect -337 -188 -303 188
rect -209 -188 -175 188
rect -81 -188 -47 188
rect 47 -188 81 188
rect 175 -188 209 188
rect 303 -188 337 188
<< metal1 >>
rect -287 281 287 287
rect -287 247 -275 281
rect 275 247 287 281
rect -287 241 287 247
rect -343 188 -297 200
rect -343 -188 -337 188
rect -303 -188 -297 188
rect -343 -200 -297 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -87 188 -41 200
rect -87 -188 -81 188
rect -47 -188 -41 188
rect -87 -200 -41 -188
rect 41 188 87 200
rect 41 -188 47 188
rect 81 -188 87 188
rect 41 -200 87 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 297 188 343 200
rect 297 -188 303 188
rect 337 -188 343 188
rect 297 -200 343 -188
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -434 -366 434 366
string parameters w 2 l 0.35 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
