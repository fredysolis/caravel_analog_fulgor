magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect -235 1684 483 1772
<< pwell >>
rect -235 1054 -139 1066
rect 409 1064 483 1066
rect -235 922 -131 1054
rect -235 556 -139 922
rect 387 556 483 1064
rect -235 468 483 556
<< psubdiff >>
rect -199 861 -165 934
rect -199 626 -165 655
rect 413 872 447 934
rect 413 626 447 666
rect -199 592 -23 626
rect 255 592 447 626
rect -31 504 -7 538
rect 255 504 279 538
<< nsubdiff >>
rect -127 1702 -103 1736
rect 351 1702 375 1736
<< psubdiffcont >>
rect -199 655 -165 861
rect 413 666 447 872
rect -7 504 255 538
<< nsubdiffcont >>
rect -103 1702 351 1736
<< poly >>
rect -35 1193 31 1217
rect -35 1111 -25 1193
rect 9 1111 31 1193
rect 253 1125 319 1259
rect -35 948 31 1111
rect 157 1059 319 1125
rect 157 1053 223 1059
rect 157 971 172 1053
rect 206 971 223 1053
rect -35 882 61 948
rect 157 878 223 971
<< polycont >>
rect -25 1111 9 1193
rect 172 971 206 1053
<< locali >>
rect -25 1193 9 1209
rect -25 1095 9 1111
rect 172 1053 206 1069
rect 172 955 206 971
rect -199 861 -165 934
rect -199 626 -165 655
rect 413 872 447 934
rect 413 626 447 666
rect -199 592 -103 626
rect 351 592 447 626
<< viali >>
rect -199 1702 -103 1736
rect -103 1702 351 1736
rect 351 1702 447 1736
rect -199 1614 447 1648
rect -25 1111 9 1193
rect 172 971 206 1053
rect -103 592 351 626
rect -103 504 -7 538
rect -7 504 255 538
rect 255 504 351 538
<< metal1 >>
rect -235 1736 483 1742
rect -235 1702 -199 1736
rect 447 1702 483 1736
rect -235 1648 483 1702
rect -235 1614 -199 1648
rect 447 1614 483 1648
rect -235 1608 483 1614
rect -91 1463 -45 1608
rect 293 1463 339 1608
rect 293 1375 329 1463
rect 101 1256 147 1297
rect 101 1210 337 1256
rect -31 1193 15 1205
rect -31 1186 -25 1193
rect -235 1120 -25 1186
rect -31 1111 -25 1120
rect 9 1111 15 1193
rect -31 1099 15 1111
rect 166 1053 212 1065
rect 166 1025 172 1053
rect -235 971 172 1025
rect 206 971 212 1053
rect -235 959 212 971
rect 291 931 337 1210
rect 101 885 337 931
rect 101 855 147 885
rect 5 632 51 774
rect 197 632 243 776
rect -235 626 483 632
rect -235 592 -103 626
rect 351 592 483 626
rect -235 538 483 592
rect -235 504 -103 538
rect 351 504 483 538
rect -235 498 483 504
use sky130_fd_pr__nfet_01v8_C3YG4M  sky130_fd_pr__nfet_01v8_C3YG4M_0
timestamp 1624049879
transform 1 0 124 0 1 811
box -263 -255 263 255
use sky130_fd_pr__pfet_01v8_4F35BC  sky130_fd_pr__pfet_01v8_4F35BC_0
timestamp 1624049879
transform 1 0 124 0 1 1375
box -359 -309 359 309
<< labels >>
rlabel metal1 -235 1648 483 1702 1 vdd
rlabel metal1 -235 538 483 592 1 vss
rlabel metal1 -235 1120 -25 1186 1 A
rlabel metal1 -235 959 172 1025 1 B
rlabel metal1 291 885 337 1256 1 out
<< end >>
