magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< pwell >>
rect -1127 -285 1127 285
<< nmos >>
rect -927 -75 -897 75
rect -831 -75 -801 75
rect -735 -75 -705 75
rect -639 -75 -609 75
rect -543 -75 -513 75
rect -447 -75 -417 75
rect -351 -75 -321 75
rect -255 -75 -225 75
rect -159 -75 -129 75
rect -63 -75 -33 75
rect 33 -75 63 75
rect 129 -75 159 75
rect 225 -75 255 75
rect 321 -75 351 75
rect 417 -75 447 75
rect 513 -75 543 75
rect 609 -75 639 75
rect 705 -75 735 75
rect 801 -75 831 75
rect 897 -75 927 75
<< ndiff >>
rect -989 63 -927 75
rect -989 -63 -977 63
rect -943 -63 -927 63
rect -989 -75 -927 -63
rect -897 63 -831 75
rect -897 -63 -881 63
rect -847 -63 -831 63
rect -897 -75 -831 -63
rect -801 63 -735 75
rect -801 -63 -785 63
rect -751 -63 -735 63
rect -801 -75 -735 -63
rect -705 63 -639 75
rect -705 -63 -689 63
rect -655 -63 -639 63
rect -705 -75 -639 -63
rect -609 63 -543 75
rect -609 -63 -593 63
rect -559 -63 -543 63
rect -609 -75 -543 -63
rect -513 63 -447 75
rect -513 -63 -497 63
rect -463 -63 -447 63
rect -513 -75 -447 -63
rect -417 63 -351 75
rect -417 -63 -401 63
rect -367 -63 -351 63
rect -417 -75 -351 -63
rect -321 63 -255 75
rect -321 -63 -305 63
rect -271 -63 -255 63
rect -321 -75 -255 -63
rect -225 63 -159 75
rect -225 -63 -209 63
rect -175 -63 -159 63
rect -225 -75 -159 -63
rect -129 63 -63 75
rect -129 -63 -113 63
rect -79 -63 -63 63
rect -129 -75 -63 -63
rect -33 63 33 75
rect -33 -63 -17 63
rect 17 -63 33 63
rect -33 -75 33 -63
rect 63 63 129 75
rect 63 -63 79 63
rect 113 -63 129 63
rect 63 -75 129 -63
rect 159 63 225 75
rect 159 -63 175 63
rect 209 -63 225 63
rect 159 -75 225 -63
rect 255 63 321 75
rect 255 -63 271 63
rect 305 -63 321 63
rect 255 -75 321 -63
rect 351 63 417 75
rect 351 -63 367 63
rect 401 -63 417 63
rect 351 -75 417 -63
rect 447 63 513 75
rect 447 -63 463 63
rect 497 -63 513 63
rect 447 -75 513 -63
rect 543 63 609 75
rect 543 -63 559 63
rect 593 -63 609 63
rect 543 -75 609 -63
rect 639 63 705 75
rect 639 -63 655 63
rect 689 -63 705 63
rect 639 -75 705 -63
rect 735 63 801 75
rect 735 -63 751 63
rect 785 -63 801 63
rect 735 -75 801 -63
rect 831 63 897 75
rect 831 -63 847 63
rect 881 -63 897 63
rect 831 -75 897 -63
rect 927 63 989 75
rect 927 -63 943 63
rect 977 -63 989 63
rect 927 -75 989 -63
<< ndiffc >>
rect -977 -63 -943 63
rect -881 -63 -847 63
rect -785 -63 -751 63
rect -689 -63 -655 63
rect -593 -63 -559 63
rect -497 -63 -463 63
rect -401 -63 -367 63
rect -305 -63 -271 63
rect -209 -63 -175 63
rect -113 -63 -79 63
rect -17 -63 17 63
rect 79 -63 113 63
rect 175 -63 209 63
rect 271 -63 305 63
rect 367 -63 401 63
rect 463 -63 497 63
rect 559 -63 593 63
rect 655 -63 689 63
rect 751 -63 785 63
rect 847 -63 881 63
rect 943 -63 977 63
<< psubdiff >>
rect -1057 -249 -995 -215
rect 995 -249 1057 -215
<< psubdiffcont >>
rect -995 -249 995 -215
<< poly >>
rect -927 97 -33 163
rect -927 75 -897 97
rect -831 75 -801 97
rect -735 75 -705 97
rect -639 75 -609 97
rect -543 75 -513 97
rect -447 75 -417 97
rect -351 75 -321 97
rect -255 75 -225 97
rect -159 75 -129 97
rect -63 75 -33 97
rect 33 97 927 163
rect 33 75 63 97
rect 129 75 159 97
rect 225 75 255 97
rect 321 75 351 97
rect 417 75 447 97
rect 513 75 543 97
rect 609 75 639 97
rect 705 75 735 97
rect 801 75 831 97
rect 897 75 927 97
rect -927 -101 -897 -75
rect -831 -101 -801 -75
rect -735 -101 -705 -75
rect -639 -101 -609 -75
rect -543 -101 -513 -75
rect -447 -101 -417 -75
rect -351 -101 -321 -75
rect -255 -101 -225 -75
rect -159 -101 -129 -75
rect -63 -101 -33 -75
rect 33 -101 63 -75
rect 129 -101 159 -75
rect 225 -101 255 -75
rect 321 -101 351 -75
rect 417 -101 447 -75
rect 513 -101 543 -75
rect 609 -101 639 -75
rect 705 -101 735 -75
rect 801 -101 831 -75
rect 897 -101 927 -75
<< locali >>
rect -977 63 -943 79
rect -977 -79 -943 -63
rect -881 63 -847 79
rect -881 -79 -847 -63
rect -785 63 -751 79
rect -785 -79 -751 -63
rect -689 63 -655 79
rect -689 -79 -655 -63
rect -593 63 -559 79
rect -593 -79 -559 -63
rect -497 63 -463 79
rect -497 -79 -463 -63
rect -401 63 -367 79
rect -401 -79 -367 -63
rect -305 63 -271 79
rect -305 -79 -271 -63
rect -209 63 -175 79
rect -209 -79 -175 -63
rect -113 63 -79 79
rect -113 -79 -79 -63
rect -17 63 17 79
rect -17 -79 17 -63
rect 79 63 113 79
rect 79 -79 113 -63
rect 175 63 209 79
rect 175 -79 209 -63
rect 271 63 305 79
rect 271 -79 305 -63
rect 367 63 401 79
rect 367 -79 401 -63
rect 463 63 497 79
rect 463 -79 497 -63
rect 559 63 593 79
rect 559 -79 593 -63
rect 655 63 689 79
rect 655 -79 689 -63
rect 751 63 785 79
rect 751 -79 785 -63
rect 847 63 881 79
rect 847 -79 881 -63
rect 943 63 977 79
rect 943 -79 977 -63
rect -1057 -249 -995 -215
rect 995 -249 1057 -215
<< viali >>
rect -977 -63 -943 63
rect -881 -63 -847 63
rect -785 -63 -751 63
rect -689 -63 -655 63
rect -593 -63 -559 63
rect -497 -63 -463 63
rect -401 -63 -367 63
rect -305 -63 -271 63
rect -209 -63 -175 63
rect -113 -63 -79 63
rect -17 -63 17 63
rect 79 -63 113 63
rect 175 -63 209 63
rect 271 -63 305 63
rect 367 -63 401 63
rect 463 -63 497 63
rect 559 -63 593 63
rect 655 -63 689 63
rect 751 -63 785 63
rect 847 -63 881 63
rect 943 -63 977 63
<< metal1 >>
rect -983 63 -937 75
rect -983 -63 -977 63
rect -943 -63 -937 63
rect -983 -75 -937 -63
rect -887 63 -841 75
rect -887 -63 -881 63
rect -847 -63 -841 63
rect -887 -75 -841 -63
rect -791 63 -745 75
rect -791 -63 -785 63
rect -751 -63 -745 63
rect -791 -75 -745 -63
rect -695 63 -649 75
rect -695 -63 -689 63
rect -655 -63 -649 63
rect -695 -75 -649 -63
rect -599 63 -553 75
rect -599 -63 -593 63
rect -559 -63 -553 63
rect -599 -75 -553 -63
rect -503 63 -457 75
rect -503 -63 -497 63
rect -463 -63 -457 63
rect -503 -75 -457 -63
rect -407 63 -361 75
rect -407 -63 -401 63
rect -367 -63 -361 63
rect -407 -75 -361 -63
rect -311 63 -265 75
rect -311 -63 -305 63
rect -271 -63 -265 63
rect -311 -75 -265 -63
rect -215 63 -169 75
rect -215 -63 -209 63
rect -175 -63 -169 63
rect -215 -75 -169 -63
rect -119 63 -73 75
rect -119 -63 -113 63
rect -79 -63 -73 63
rect -119 -75 -73 -63
rect -23 63 23 75
rect -23 -63 -17 63
rect 17 -63 23 63
rect -23 -75 23 -63
rect 73 63 119 75
rect 73 -63 79 63
rect 113 -63 119 63
rect 73 -75 119 -63
rect 169 63 215 75
rect 169 -63 175 63
rect 209 -63 215 63
rect 169 -75 215 -63
rect 265 63 311 75
rect 265 -63 271 63
rect 305 -63 311 63
rect 265 -75 311 -63
rect 361 63 407 75
rect 361 -63 367 63
rect 401 -63 407 63
rect 361 -75 407 -63
rect 457 63 503 75
rect 457 -63 463 63
rect 497 -63 503 63
rect 457 -75 503 -63
rect 553 63 599 75
rect 553 -63 559 63
rect 593 -63 599 63
rect 553 -75 599 -63
rect 649 63 695 75
rect 649 -63 655 63
rect 689 -63 695 63
rect 649 -75 695 -63
rect 745 63 791 75
rect 745 -63 751 63
rect 785 -63 791 63
rect 745 -75 791 -63
rect 841 63 887 75
rect 841 -63 847 63
rect 881 -63 887 63
rect 841 -75 887 -63
rect 937 63 983 75
rect 937 -63 943 63
rect 977 -63 983 63
rect 937 -75 983 -63
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1074 -232 1074 232
string parameters w 0.75 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
