magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< pwell >>
rect -311 -335 311 335
<< nmos >>
rect -111 -125 -81 125
rect -15 -125 15 125
rect 81 -125 111 125
<< ndiff >>
rect -173 113 -111 125
rect -173 -113 -161 113
rect -127 -113 -111 113
rect -173 -125 -111 -113
rect -81 113 -15 125
rect -81 -113 -65 113
rect -31 -113 -15 113
rect -81 -125 -15 -113
rect 15 113 81 125
rect 15 -113 31 113
rect 65 -113 81 113
rect 15 -125 81 -113
rect 111 113 173 125
rect 111 -113 127 113
rect 161 -113 173 113
rect 111 -125 173 -113
<< ndiffc >>
rect -161 -113 -127 113
rect -65 -113 -31 113
rect 31 -113 65 113
rect 127 -113 161 113
<< psubdiff >>
rect -275 203 -241 265
rect 241 203 275 265
rect -275 -265 -241 -203
rect 241 -265 275 -203
rect -275 -299 -179 -265
rect 179 -299 275 -265
<< psubdiffcont >>
rect -275 -203 -241 203
rect 241 -203 275 203
rect -179 -299 179 -265
<< poly >>
rect -111 125 -81 151
rect -15 125 15 151
rect 81 125 111 151
rect -111 -151 -81 -125
rect -15 -151 15 -125
rect 81 -151 111 -125
<< locali >>
rect -275 203 -241 265
rect 241 203 275 265
rect -161 113 -127 129
rect -161 -129 -127 -113
rect -65 113 -31 129
rect -65 -129 -31 -113
rect 31 113 65 129
rect 31 -129 65 -113
rect 127 113 161 129
rect 127 -129 161 -113
rect -275 -265 -241 -203
rect 241 -265 275 -203
rect -275 -299 -179 -265
rect 179 -299 275 -265
<< viali >>
rect -161 -113 -127 113
rect -65 -113 -31 113
rect 31 -113 65 113
rect 127 -113 161 113
<< metal1 >>
rect -167 113 -121 125
rect -167 -113 -161 113
rect -127 -113 -121 113
rect -167 -125 -121 -113
rect -71 113 -25 125
rect -71 -113 -65 113
rect -31 -113 -25 113
rect -71 -125 -25 -113
rect 25 113 71 125
rect 25 -113 31 113
rect 65 -113 71 113
rect 25 -125 71 -113
rect 121 113 167 125
rect 121 -113 127 113
rect 161 -113 167 113
rect 121 -125 167 -113
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -258 -282 258 282
string parameters w 1.25 l 0.150 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
