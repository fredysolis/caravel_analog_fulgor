magic
tech sky130A
magscale 1 2
timestamp 1624885207
<< nwell >>
rect 559 2292 1181 3068
rect 559 0 1181 776
<< pwell >>
rect 559 1729 1740 2292
rect 460 1400 1740 1729
rect 559 776 1740 1400
<< psubdiff >>
rect 433 2222 654 2256
rect 489 1718 1242 1752
rect 487 1316 1249 1350
rect 1000 812 1307 846
<< poly >>
rect 741 2104 1000 2170
rect 740 898 999 964
<< locali >>
rect 433 2222 462 2256
rect 556 2222 654 2256
rect 483 1718 1265 1752
rect 489 1316 1256 1350
rect 1028 812 1205 846
rect 1299 812 1310 846
<< viali >>
rect 462 2222 556 2256
rect 1205 812 1299 846
<< metal1 >>
rect 523 3027 1200 3038
rect 523 2998 1253 3027
rect -1244 2944 1740 2998
rect 523 2940 1195 2944
rect 523 2904 1198 2940
rect -131 2240 -121 2344
rect 450 2256 596 2262
rect 450 2222 462 2256
rect 556 2222 596 2256
rect 450 2216 596 2222
rect 219 1802 229 1854
rect 361 1814 371 1854
rect 361 1802 373 1814
rect 1393 1811 1403 1863
rect 1486 1811 1496 1863
rect 587 1712 636 1758
rect -1244 1498 69 1570
rect 1105 1310 1167 1356
rect 219 1254 231 1266
rect 221 1214 231 1254
rect 361 1254 373 1266
rect 361 1214 371 1254
rect 1392 1208 1402 1260
rect 1486 1208 1496 1260
rect 1157 846 1311 852
rect -91 724 -81 828
rect 1157 812 1205 846
rect 1299 812 1311 846
rect 1157 806 1311 812
rect 559 124 1181 164
rect -1244 70 1740 124
rect 559 30 1181 70
<< via1 >>
rect -190 2240 -131 2344
rect 229 1802 361 1854
rect 1403 1811 1486 1863
rect 231 1214 361 1266
rect 1402 1208 1486 1260
rect -150 724 -91 828
<< metal2 >>
rect -190 2344 -131 2354
rect -131 2266 40 2318
rect -190 2230 -131 2240
rect -12 1854 40 2266
rect 1521 2258 1577 2369
rect 229 1854 361 1864
rect -12 1802 229 1854
rect 229 1792 361 1802
rect 1403 1863 1486 1873
rect 1403 1801 1486 1811
rect 373 1748 429 1758
rect 1413 1722 1473 1801
rect 429 1662 1473 1722
rect 373 1626 429 1636
rect 163 1432 219 1442
rect 219 1346 1473 1406
rect 163 1310 219 1320
rect 231 1266 361 1276
rect 1413 1270 1473 1346
rect -12 1214 231 1266
rect -150 828 -91 838
rect -12 802 40 1214
rect 231 1204 361 1214
rect 1402 1260 1486 1270
rect 1402 1198 1486 1208
rect -91 750 40 802
rect -150 714 -91 724
rect 1311 699 1367 810
<< via2 >>
rect 373 1636 429 1748
rect 163 1320 219 1432
<< metal3 >>
rect -997 804 -937 2264
rect 363 1748 439 1753
rect 363 1636 373 1748
rect 429 1636 439 1748
rect 363 1631 439 1636
rect 153 1432 229 1437
rect 153 1320 163 1432
rect 219 1320 229 1432
rect 153 1315 229 1320
use clock_inverter  clock_inverter_0
timestamp 1624885207
transform 1 0 -1244 0 1 0
box 0 0 1244 3068
use latch_diff  latch_diff_1
timestamp 1624049879
transform -1 0 1707 0 -1 2352
box -33 -716 1147 2352
use latch_diff  latch_diff_0
timestamp 1624049879
transform 1 0 33 0 1 716
box -33 -716 1147 2352
<< labels >>
rlabel metal1 -1244 1498 69 1570 1 vss
rlabel metal1 -1244 2944 1740 2998 1 vdd
rlabel metal3 -997 1498 -937 1570 1 D
rlabel poly 740 898 999 964 1 CLK
rlabel poly 741 2104 1000 2170 1 nCLK
rlabel metal2 1311 699 1367 810 1 nQ
rlabel metal2 1521 2258 1577 2369 1 Q
<< end >>
