magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< viali >>
rect 126 34 1358 84
<< metal1 >>
rect 144 5172 1336 5636
rect 148 158 1340 622
rect 114 84 1370 90
rect 114 34 126 84
rect 1358 34 1370 84
rect 114 28 1370 34
use sky130_fd_pr__res_high_po_5p73_X44RQA *sky130_fd_pr__res_high_po_5p73_X44RQA_0
timestamp 1624049879
transform 1 0 739 0 1 2890
box -739 -2890 739 2890
<< labels >>
rlabel metal1 144 5172 1336 5636 1 in
rlabel viali 126 34 1358 84 1 vss
rlabel metal1 148 158 1340 622 1 out
<< end >>
