magic
tech sky130A
magscale 1 2
timestamp 1624113565
<< nwell >>
rect -51 1207 3503 1296
rect 3391 641 3503 1207
rect 3385 573 3503 641
rect 3321 -129 3503 573
rect 1777 -199 3247 -129
rect 3315 -199 3503 -129
<< pwell >>
rect -15 -103 1601 -69
<< psubdiff >>
rect -15 -103 81 -69
rect 727 -103 885 -69
rect 1531 -103 1601 -69
<< nsubdiff >>
rect -15 1226 81 1260
rect 1591 1226 1749 1260
rect 3259 1226 3355 1260
rect 3414 1075 3448 1171
rect 3414 605 3448 701
rect 3414 436 3448 533
rect 3414 -163 3448 -66
<< psubdiffcont >>
rect 81 -103 727 -69
rect 885 -103 1531 -69
<< nsubdiffcont >>
rect 81 1226 1591 1260
rect 1749 1226 3259 1260
rect 3414 701 3448 1075
rect 3414 -66 3448 436
<< viali >>
rect -15 1226 81 1260
rect 81 1226 1591 1260
rect 1591 1226 1749 1260
rect 1749 1226 3259 1260
rect 3259 1226 3355 1260
rect -15 1137 3355 1171
rect 3321 605 3355 1137
rect 3414 1075 3448 1171
rect 3414 701 3448 1075
rect 3414 605 3448 701
rect -15 -15 1601 19
rect -15 -103 81 -69
rect 81 -103 727 -69
rect 727 -103 885 -69
rect 885 -103 1531 -69
rect 1531 -103 1601 -69
rect 3321 -129 3355 533
rect 3414 436 3448 533
rect 3414 -66 3448 436
rect 3414 -163 3448 -66
<< metal1 >>
rect -51 1260 3503 1296
rect -51 1226 -15 1260
rect 3355 1226 3503 1260
rect -51 1171 3503 1226
rect -51 1137 -15 1171
rect -27 1131 3321 1137
rect 93 967 139 1131
rect 285 981 331 1131
rect 477 984 523 1131
rect 669 983 715 1131
rect 861 984 907 1131
rect 1053 982 1099 1131
rect 1245 983 1291 1131
rect 1437 984 1483 1131
rect 1761 982 1807 1131
rect 189 828 235 910
rect 381 828 427 913
rect 573 828 619 912
rect 765 828 811 909
rect 957 828 1003 912
rect 1149 828 1195 911
rect 1341 828 1387 908
rect 1533 828 1579 878
rect 189 757 235 808
rect 381 757 427 810
rect 573 757 619 811
rect 765 757 811 810
rect 957 757 1003 812
rect 1149 757 1195 810
rect 1341 757 1387 810
rect 1533 757 1579 805
rect 1837 788 1847 988
rect 1913 788 1923 988
rect 1953 981 1999 1131
rect 2029 788 2039 988
rect 2105 788 2115 988
rect 2145 982 2191 1131
rect 2221 788 2231 988
rect 2297 788 2307 988
rect 2337 987 2383 1131
rect 2413 788 2423 988
rect 2489 788 2499 988
rect 2529 983 2575 1131
rect 2605 788 2615 988
rect 2681 788 2691 988
rect 2721 983 2767 1131
rect 2797 788 2807 988
rect 2873 788 2883 988
rect 2913 982 2959 1131
rect 2989 788 2999 988
rect 3065 788 3075 988
rect 3105 982 3151 1131
rect 3181 788 3191 988
rect 3257 788 3267 988
rect 131 747 1579 757
rect 131 726 3205 747
rect 121 658 131 726
rect 1541 658 3205 726
rect 3315 605 3321 1131
rect 3355 605 3414 1171
rect 3448 605 3503 1171
rect 3315 533 3503 605
rect 137 393 1477 499
rect 189 329 235 393
rect 381 335 427 393
rect 573 343 619 393
rect 659 391 952 393
rect 1973 390 3195 446
rect 93 25 139 177
rect 285 25 331 185
rect 477 25 523 190
rect 669 25 715 188
rect 897 25 943 185
rect 973 159 983 359
rect 1049 159 1059 359
rect 1089 25 1135 188
rect 1165 159 1175 359
rect 1241 159 1251 359
rect 1281 25 1327 188
rect 1357 159 1367 359
rect 1433 159 1443 359
rect 1473 25 1519 187
rect -27 19 1777 25
rect -51 -15 -15 19
rect 1601 -15 1777 19
rect -51 -69 1777 -15
rect -51 -103 -15 -69
rect 1601 -103 1777 -69
rect -51 -123 1777 -103
rect 1921 -123 1967 -11
rect 2033 -51 2043 349
rect 2101 -51 2111 349
rect 2177 -123 2223 1
rect 2289 -51 2299 349
rect 2357 -51 2367 349
rect 2433 -123 2479 4
rect 2545 -51 2555 349
rect 2613 -51 2623 349
rect 2689 -123 2735 9
rect 2801 -51 2811 349
rect 2869 -51 2879 349
rect 2945 -123 2991 13
rect 3057 -51 3067 349
rect 3125 -51 3135 349
rect 3201 -123 3247 8
rect -51 -311 3247 -123
rect 3315 -129 3321 533
rect 3355 -129 3414 533
rect 3315 -163 3414 -129
rect 3448 -163 3503 533
rect 3315 -199 3503 -163
<< via1 >>
rect 1847 788 1913 988
rect 2039 788 2105 988
rect 2231 788 2297 988
rect 2423 788 2489 988
rect 2615 788 2681 988
rect 2807 788 2873 988
rect 2999 788 3065 988
rect 3191 788 3257 988
rect 131 658 1541 726
rect 983 159 1049 359
rect 1175 159 1241 359
rect 1367 159 1433 359
rect 2043 -51 2101 349
rect 2299 -51 2357 349
rect 2555 -51 2613 349
rect 2811 -51 2869 349
rect 3067 -51 3125 349
<< metal2 >>
rect 1847 988 3257 998
rect 1913 788 2039 988
rect 2105 788 2231 988
rect 2297 788 2423 988
rect 2489 788 2615 988
rect 2681 788 2807 988
rect 2873 788 2999 988
rect 3065 788 3191 988
rect 1847 778 3257 788
rect 131 726 1541 736
rect 131 648 1541 658
rect 990 369 1423 648
rect 983 359 1433 369
rect 1049 159 1175 359
rect 1241 159 1367 359
rect 983 149 1433 159
rect 2043 349 3125 778
rect 2101 -51 2299 349
rect 2357 -51 2555 349
rect 2613 -51 2811 349
rect 2869 -51 3067 349
rect 2043 -61 3125 -51
use sky130_fd_pr__pfet_01v8_VCU74W  sky130_fd_pr__pfet_01v8_VCU74W_0
timestamp 1623969746
transform 1 0 836 0 1 888
box -887 -319 887 319
use sky130_fd_pr__pfet_01v8_VCU74W  sky130_fd_pr__pfet_01v8_VCU74W_1
timestamp 1623969746
transform 1 0 2504 0 1 888
box -887 -319 887 319
use sky130_fd_pr__pfet_01v8_lvt_D3F744  sky130_fd_pr__pfet_01v8_lvt_D3F744_0
timestamp 1623976832
transform 1 0 2584 0 1 185
box -807 -384 807 384
use sky130_fd_pr__nfet_01v8_lvt_9B2JY7  sky130_fd_pr__nfet_01v8_lvt_9B2JY7_0 
timestamp 1624020979
transform 1 0 404 0 1 259
box -455 -310 455 310
use sky130_fd_pr__nfet_01v8_lvt_9B2JY7  sky130_fd_pr__nfet_01v8_lvt_9B2JY7_1
timestamp 1624020979
transform 1 0 1208 0 1 259
box -455 -310 455 310
<< labels >>
rlabel metal2 3060 554 3092 593 1 out
rlabel metal1 195 395 227 434 1 iref
rlabel metal1 -18 -180 14 -141 1 avss1p8
rlabel metal1 -9 1181 23 1220 1 avdd1p8
rlabel metal1 1973 390 3195 446 1 in
<< end >>
