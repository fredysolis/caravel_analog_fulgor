magic
tech sky130A
magscale 1 2
timestamp 1624020979
<< pwell >>
rect -455 188 455 310
rect -455 122 -205 188
rect -203 122 -15 188
rect -12 122 178 188
rect 180 122 455 188
rect -455 -310 455 122
<< nmoslvt >>
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
<< ndiff >>
rect -317 88 -255 100
rect -317 -88 -305 88
rect -271 -88 -255 88
rect -317 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 317 100
rect 255 -88 271 88
rect 305 -88 317 88
rect 255 -100 317 -88
<< ndiffc >>
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
<< psubdiff >>
rect -419 240 -323 274
rect 323 240 419 274
rect -419 178 -385 240
rect 385 178 419 240
rect -419 -240 -385 -178
rect 385 -240 419 -178
rect -419 -274 -323 -240
rect 323 -274 419 -240
<< psubdiffcont >>
rect -323 240 323 274
rect -419 -178 -385 178
rect 385 -178 419 178
rect -323 -274 323 -240
<< poly >>
rect -271 172 273 188
rect -271 138 -255 172
rect -221 138 -161 172
rect -127 138 -65 172
rect -31 138 31 172
rect 65 138 128 172
rect 162 138 223 172
rect 257 138 273 172
rect -271 122 273 138
rect -255 100 -225 122
rect -159 100 -129 122
rect -63 100 -33 122
rect 33 100 63 122
rect 129 100 159 122
rect 225 100 255 122
rect -255 -126 -225 -100
rect -159 -126 -129 -100
rect -63 -126 -33 -100
rect 33 -126 63 -100
rect 129 -126 159 -100
rect 225 -126 255 -100
<< polycont >>
rect -255 138 -221 172
rect -161 138 -127 172
rect -65 138 -31 172
rect 31 138 65 172
rect 128 138 162 172
rect 223 138 257 172
<< locali >>
rect -419 240 -323 274
rect 323 240 419 274
rect -419 178 -385 240
rect 385 178 419 240
rect -271 138 -255 172
rect 257 138 273 172
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect -419 -240 -385 -178
rect 385 -240 419 -178
rect -419 -274 -323 -240
rect 323 -274 419 -240
<< viali >>
rect -255 138 -221 172
rect -221 138 -161 172
rect -161 138 -127 172
rect -127 138 -65 172
rect -65 138 -31 172
rect -31 138 31 172
rect 31 138 65 172
rect 65 138 128 172
rect 128 138 162 172
rect 162 138 223 172
rect 223 138 257 172
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
<< metal1 >>
rect -267 172 269 178
rect -267 138 -255 172
rect 257 138 269 172
rect -267 132 269 138
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -402 -257 402 257
string parameters w 1 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
