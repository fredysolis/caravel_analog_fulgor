magic
tech sky130A
magscale 1 2
timestamp 1624018159
<< error_p >>
rect -2890 8140 -2770 13200
rect -4483 8000 -2770 8140
rect -2650 8140 -2530 13200
rect 2429 8140 2549 13200
rect -2650 8000 2549 8140
rect 2669 8140 2789 13200
rect 7748 8140 7868 13200
rect 2669 8000 7868 8140
rect 7988 8140 8108 13200
rect 7988 8000 13287 8140
rect -4483 7760 -2770 7900
rect -2890 2840 -2770 7760
rect -4483 2700 -2770 2840
rect -2650 7760 2549 7900
rect -2650 2840 -2530 7760
rect 2429 2840 2549 7760
rect -2650 2700 2549 2840
rect 2669 7760 7868 7900
rect 2669 2840 2789 7760
rect 7748 2840 7868 7760
rect 2669 2700 7868 2840
rect 7988 7760 13287 7900
rect 7988 2840 8108 7760
rect 7988 2700 13287 2840
rect -4483 2460 -2770 2600
rect -2890 -2460 -2770 2460
rect -4483 -2600 -2770 -2460
rect -2650 2460 2549 2600
rect -2650 -2460 -2530 2460
rect 2429 -2460 2549 2460
rect -2650 -2600 2549 -2460
rect 2669 2460 7868 2600
rect 2669 -2460 2789 2460
rect 7748 -2460 7868 2460
rect 2669 -2600 7868 -2460
rect 7988 2460 13287 2600
rect 7988 -2460 8108 2460
rect 7988 -2600 13287 -2460
rect -4483 -2840 -2770 -2700
rect -2890 -7760 -2770 -2840
rect -4483 -7900 -2770 -7760
rect -2650 -2840 2549 -2700
rect -2650 -7760 -2530 -2840
rect 2429 -7760 2549 -2840
rect -2650 -7900 2549 -7760
rect 2669 -2840 7868 -2700
rect 2669 -7760 2789 -2840
rect 7748 -7760 7868 -2840
rect 2669 -7900 7868 -7760
rect 7988 -2840 13287 -2700
rect 7988 -7760 8108 -2840
rect 7988 -7900 13287 -7760
rect -4483 -8140 -2770 -8000
rect -2890 -12071 -2770 -8140
rect -2650 -8140 2549 -8000
rect -2650 -12071 -2530 -8140
rect 2429 -12071 2549 -8140
rect 2669 -8140 7868 -8000
rect 2669 -12071 2789 -8140
rect 7748 -12071 7868 -8140
rect 7988 -8140 13287 -8000
rect 7988 -12071 8108 -8140
<< metal3 >>
rect -13288 8000 -8089 13200
rect -7969 8000 -2770 13200
rect -2650 8000 2549 13200
rect 2669 8000 7868 13200
rect 7988 13172 13287 13200
rect 7988 8028 13203 13172
rect 13267 8028 13287 13172
rect 7988 8000 13287 8028
rect -13288 2700 -8089 7900
rect -7969 2700 -2770 7900
rect -2650 2700 2549 7900
rect 2669 2700 7868 7900
rect 7988 7872 13287 7900
rect 7988 2728 13203 7872
rect 13267 2728 13287 7872
rect 7988 2700 13287 2728
rect -13288 -2600 -8089 2600
rect -7969 -2600 -2770 2600
rect -2650 -2600 2549 2600
rect 2669 -2600 7868 2600
rect 7988 2572 13287 2600
rect 7988 -2572 13203 2572
rect 13267 -2572 13287 2572
rect 7988 -2600 13287 -2572
rect -13288 -7900 -8089 -2700
rect -7969 -7900 -2770 -2700
rect -2650 -7900 2549 -2700
rect 2669 -7900 7868 -2700
rect 7988 -2728 13287 -2700
rect 7988 -7872 13203 -2728
rect 13267 -7872 13287 -2728
rect 7988 -7900 13287 -7872
rect -13288 -13200 -8089 -8000
rect -7969 -13200 -2770 -8000
rect -2650 -13200 2549 -8000
rect 2669 -13200 7868 -8000
rect 7988 -8028 13287 -8000
rect 7988 -13172 13203 -8028
rect 13267 -13172 13287 -8028
rect 7988 -13200 13287 -13172
<< via3 >>
rect 13203 8028 13267 13172
rect 13203 2728 13267 7872
rect 13203 -2572 13267 2572
rect 13203 -7872 13267 -2728
rect 13203 -13172 13267 -8028
<< mimcap >>
rect -13188 13060 -8188 13100
rect -13188 8140 -13148 13060
rect -8228 8140 -8188 13060
rect -13188 8100 -8188 8140
rect -7869 13060 -2869 13100
rect -7869 8140 -7829 13060
rect -2909 8140 -2869 13060
rect -7869 8100 -2869 8140
rect -2550 13060 2450 13100
rect -2550 8140 -2510 13060
rect 2410 8140 2450 13060
rect -2550 8100 2450 8140
rect 2769 13060 7769 13100
rect 2769 8140 2809 13060
rect 7729 8140 7769 13060
rect 2769 8100 7769 8140
rect 8088 13060 13088 13100
rect 8088 8140 8128 13060
rect 13048 8140 13088 13060
rect 8088 8100 13088 8140
rect -13188 7760 -8188 7800
rect -13188 2840 -13148 7760
rect -8228 2840 -8188 7760
rect -13188 2800 -8188 2840
rect -7869 7760 -2869 7800
rect -7869 2840 -7829 7760
rect -2909 2840 -2869 7760
rect -7869 2800 -2869 2840
rect -2550 7760 2450 7800
rect -2550 2840 -2510 7760
rect 2410 2840 2450 7760
rect -2550 2800 2450 2840
rect 2769 7760 7769 7800
rect 2769 2840 2809 7760
rect 7729 2840 7769 7760
rect 2769 2800 7769 2840
rect 8088 7760 13088 7800
rect 8088 2840 8128 7760
rect 13048 2840 13088 7760
rect 8088 2800 13088 2840
rect -13188 2460 -8188 2500
rect -13188 -2460 -13148 2460
rect -8228 -2460 -8188 2460
rect -13188 -2500 -8188 -2460
rect -7869 2460 -2869 2500
rect -7869 -2460 -7829 2460
rect -2909 -2460 -2869 2460
rect -7869 -2500 -2869 -2460
rect -2550 2460 2450 2500
rect -2550 -2460 -2510 2460
rect 2410 -2460 2450 2460
rect -2550 -2500 2450 -2460
rect 2769 2460 7769 2500
rect 2769 -2460 2809 2460
rect 7729 -2460 7769 2460
rect 2769 -2500 7769 -2460
rect 8088 2460 13088 2500
rect 8088 -2460 8128 2460
rect 13048 -2460 13088 2460
rect 8088 -2500 13088 -2460
rect -13188 -2840 -8188 -2800
rect -13188 -7760 -13148 -2840
rect -8228 -7760 -8188 -2840
rect -13188 -7800 -8188 -7760
rect -7869 -2840 -2869 -2800
rect -7869 -7760 -7829 -2840
rect -2909 -7760 -2869 -2840
rect -7869 -7800 -2869 -7760
rect -2550 -2840 2450 -2800
rect -2550 -7760 -2510 -2840
rect 2410 -7760 2450 -2840
rect -2550 -7800 2450 -7760
rect 2769 -2840 7769 -2800
rect 2769 -7760 2809 -2840
rect 7729 -7760 7769 -2840
rect 2769 -7800 7769 -7760
rect 8088 -2840 13088 -2800
rect 8088 -7760 8128 -2840
rect 13048 -7760 13088 -2840
rect 8088 -7800 13088 -7760
rect -13188 -8140 -8188 -8100
rect -13188 -13060 -13148 -8140
rect -8228 -13060 -8188 -8140
rect -13188 -13100 -8188 -13060
rect -7869 -8140 -2869 -8100
rect -7869 -13060 -7829 -8140
rect -2909 -13060 -2869 -8140
rect -7869 -13100 -2869 -13060
rect -2550 -8140 2450 -8100
rect -2550 -13060 -2510 -8140
rect 2410 -13060 2450 -8140
rect -2550 -13100 2450 -13060
rect 2769 -8140 7769 -8100
rect 2769 -13060 2809 -8140
rect 7729 -13060 7769 -8140
rect 2769 -13100 7769 -13060
rect 8088 -8140 13088 -8100
rect 8088 -13060 8128 -8140
rect 13048 -13060 13088 -8140
rect 8088 -13100 13088 -13060
<< mimcapcontact >>
rect -13148 8140 -8228 13060
rect -7829 8140 -2909 13060
rect -2510 8140 2410 13060
rect 2809 8140 7729 13060
rect 8128 8140 13048 13060
rect -13148 2840 -8228 7760
rect -7829 2840 -2909 7760
rect -2510 2840 2410 7760
rect 2809 2840 7729 7760
rect 8128 2840 13048 7760
rect -13148 -2460 -8228 2460
rect -7829 -2460 -2909 2460
rect -2510 -2460 2410 2460
rect 2809 -2460 7729 2460
rect 8128 -2460 13048 2460
rect -13148 -7760 -8228 -2840
rect -7829 -7760 -2909 -2840
rect -2510 -7760 2410 -2840
rect 2809 -7760 7729 -2840
rect 8128 -7760 13048 -2840
rect -13148 -13060 -8228 -8140
rect -7829 -13060 -2909 -8140
rect -2510 -13060 2410 -8140
rect 2809 -13060 7729 -8140
rect 8128 -13060 13048 -8140
<< metal4 >>
rect 13187 13172 13283 13188
rect -13149 13060 -8227 13061
rect -13149 8140 -13148 13060
rect -8228 11100 -8227 13060
rect -7830 13060 -2908 13061
rect -7830 11100 -7829 13060
rect -8228 10100 -7829 11100
rect -8228 8140 -8227 10100
rect -13149 8139 -8227 8140
rect -7830 8140 -7829 10100
rect -2909 11100 -2908 13060
rect -2511 13060 2411 13061
rect -2511 11100 -2510 13060
rect -2909 10100 -2510 11100
rect -2909 8140 -2908 10100
rect -7830 8139 -2908 8140
rect -2511 8140 -2510 10100
rect 2410 11100 2411 13060
rect 2808 13060 7730 13061
rect 2808 11100 2809 13060
rect 2410 10100 2809 11100
rect 2410 8140 2411 10100
rect -2511 8139 2411 8140
rect 2808 8140 2809 10100
rect 7729 11100 7730 13060
rect 8127 13060 13049 13061
rect 8127 11100 8128 13060
rect 7729 10100 8128 11100
rect 7729 8140 7730 10100
rect 2808 8139 7730 8140
rect 8127 8140 8128 10100
rect 13048 8140 13049 13060
rect 8127 8139 13049 8140
rect -11188 7761 -10188 8139
rect -5869 7761 -4869 8139
rect -551 7761 449 8139
rect 4767 7761 5767 8139
rect 10085 7761 11085 8139
rect 13187 8028 13203 13172
rect 13267 8028 13283 13172
rect 13187 8012 13283 8028
rect 13187 7872 13283 7888
rect -13149 7760 -8227 7761
rect -13149 2840 -13148 7760
rect -8228 5800 -8227 7760
rect -7830 7760 -2908 7761
rect -7830 5800 -7829 7760
rect -8228 4800 -7829 5800
rect -8228 2840 -8227 4800
rect -13149 2839 -8227 2840
rect -7830 2840 -7829 4800
rect -2909 5800 -2908 7760
rect -2511 7760 2411 7761
rect -2511 5800 -2510 7760
rect -2909 4800 -2510 5800
rect -2909 2840 -2908 4800
rect -7830 2839 -2908 2840
rect -2511 2840 -2510 4800
rect 2410 5800 2411 7760
rect 2808 7760 7730 7761
rect 2808 5800 2809 7760
rect 2410 4800 2809 5800
rect 2410 2840 2411 4800
rect -2511 2839 2411 2840
rect 2808 2840 2809 4800
rect 7729 5800 7730 7760
rect 8127 7760 13049 7761
rect 8127 5800 8128 7760
rect 7729 4800 8128 5800
rect 7729 2840 7730 4800
rect 2808 2839 7730 2840
rect 8127 2840 8128 4800
rect 13048 2840 13049 7760
rect 8127 2839 13049 2840
rect -11188 2461 -10188 2839
rect -5869 2461 -4869 2839
rect -551 2461 449 2839
rect 4767 2461 5767 2839
rect 10085 2461 11085 2839
rect 13187 2728 13203 7872
rect 13267 2728 13283 7872
rect 13187 2712 13283 2728
rect 13187 2572 13283 2588
rect -13149 2460 -8227 2461
rect -13149 -2460 -13148 2460
rect -8228 500 -8227 2460
rect -7830 2460 -2908 2461
rect -7830 500 -7829 2460
rect -8228 -500 -7829 500
rect -8228 -2460 -8227 -500
rect -13149 -2461 -8227 -2460
rect -7830 -2460 -7829 -500
rect -2909 500 -2908 2460
rect -2511 2460 2411 2461
rect -2511 500 -2510 2460
rect -2909 -500 -2510 500
rect -2909 -2460 -2908 -500
rect -7830 -2461 -2908 -2460
rect -2511 -2460 -2510 -500
rect 2410 500 2411 2460
rect 2808 2460 7730 2461
rect 2808 500 2809 2460
rect 2410 -500 2809 500
rect 2410 -2460 2411 -500
rect -2511 -2461 2411 -2460
rect 2808 -2460 2809 -500
rect 7729 500 7730 2460
rect 8127 2460 13049 2461
rect 8127 500 8128 2460
rect 7729 -500 8128 500
rect 7729 -2460 7730 -500
rect 2808 -2461 7730 -2460
rect 8127 -2460 8128 -500
rect 13048 -2460 13049 2460
rect 8127 -2461 13049 -2460
rect -11188 -2839 -10188 -2461
rect -5869 -2839 -4869 -2461
rect -551 -2839 449 -2461
rect 4767 -2839 5767 -2461
rect 10085 -2839 11085 -2461
rect 13187 -2572 13203 2572
rect 13267 -2572 13283 2572
rect 13187 -2588 13283 -2572
rect 13187 -2728 13283 -2712
rect -13149 -2840 -8227 -2839
rect -13149 -7760 -13148 -2840
rect -8228 -4800 -8227 -2840
rect -7830 -2840 -2908 -2839
rect -7830 -4800 -7829 -2840
rect -8228 -5800 -7829 -4800
rect -8228 -7760 -8227 -5800
rect -13149 -7761 -8227 -7760
rect -7830 -7760 -7829 -5800
rect -2909 -4800 -2908 -2840
rect -2511 -2840 2411 -2839
rect -2511 -4800 -2510 -2840
rect -2909 -5800 -2510 -4800
rect -2909 -7760 -2908 -5800
rect -7830 -7761 -2908 -7760
rect -2511 -7760 -2510 -5800
rect 2410 -4800 2411 -2840
rect 2808 -2840 7730 -2839
rect 2808 -4800 2809 -2840
rect 2410 -5800 2809 -4800
rect 2410 -7760 2411 -5800
rect -2511 -7761 2411 -7760
rect 2808 -7760 2809 -5800
rect 7729 -4800 7730 -2840
rect 8127 -2840 13049 -2839
rect 8127 -4800 8128 -2840
rect 7729 -5800 8128 -4800
rect 7729 -7760 7730 -5800
rect 2808 -7761 7730 -7760
rect 8127 -7760 8128 -5800
rect 13048 -7760 13049 -2840
rect 8127 -7761 13049 -7760
rect -11188 -8139 -10188 -7761
rect -5869 -8139 -4869 -7761
rect -551 -8139 449 -7761
rect 4767 -8139 5767 -7761
rect 10085 -8139 11085 -7761
rect 13187 -7872 13203 -2728
rect 13267 -7872 13283 -2728
rect 13187 -7888 13283 -7872
rect 13187 -8028 13283 -8012
rect -13149 -8140 -8227 -8139
rect -13149 -13060 -13148 -8140
rect -8228 -10100 -8227 -8140
rect -7830 -8140 -2908 -8139
rect -7830 -10100 -7829 -8140
rect -8228 -11100 -7829 -10100
rect -8228 -13060 -8227 -11100
rect -13149 -13061 -8227 -13060
rect -7830 -13060 -7829 -11100
rect -2909 -10100 -2908 -8140
rect -2511 -8140 2411 -8139
rect -2511 -10100 -2510 -8140
rect -2909 -11100 -2510 -10100
rect -2909 -13060 -2908 -11100
rect -7830 -13061 -2908 -13060
rect -2511 -13060 -2510 -11100
rect 2410 -10100 2411 -8140
rect 2808 -8140 7730 -8139
rect 2808 -10100 2809 -8140
rect 2410 -11100 2809 -10100
rect 2410 -13060 2411 -11100
rect -2511 -13061 2411 -13060
rect 2808 -13060 2809 -11100
rect 7729 -10100 7730 -8140
rect 8127 -8140 13049 -8139
rect 8127 -10100 8128 -8140
rect 7729 -11100 8128 -10100
rect 7729 -13060 7730 -11100
rect 2808 -13061 7730 -13060
rect 8127 -13060 8128 -11100
rect 13048 -13060 13049 -8140
rect 8127 -13061 13049 -13060
rect 13187 -13172 13203 -8028
rect 13267 -13172 13283 -8028
rect 13187 -13188 13283 -13172
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 7988 8000 13188 13200
string parameters w 25 l 25 val 1.269k carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>
