magic
tech sky130A
magscale 1 2
timestamp 1623863898
<< nwell >>
rect -2017 76 2017 1196
rect -2018 -202 2017 76
rect -2017 -1367 2017 -202
<< pmoslvt >>
rect -1821 47 -1731 947
rect -1673 47 -1583 947
rect -1525 47 -1435 947
rect -1377 47 -1287 947
rect -1229 47 -1139 947
rect -1081 47 -991 947
rect -933 47 -843 947
rect -785 47 -695 947
rect -637 47 -547 947
rect -489 47 -399 947
rect -341 47 -251 947
rect -193 47 -103 947
rect -45 47 45 947
rect 103 47 193 947
rect 251 47 341 947
rect 399 47 489 947
rect 547 47 637 947
rect 695 47 785 947
rect 843 47 933 947
rect 991 47 1081 947
rect 1139 47 1229 947
rect 1287 47 1377 947
rect 1435 47 1525 947
rect 1583 47 1673 947
rect 1731 47 1821 947
rect -1821 -1219 -1731 -319
rect -1673 -1219 -1583 -319
rect -1525 -1219 -1435 -319
rect -1377 -1219 -1287 -319
rect -1229 -1219 -1139 -319
rect -1081 -1219 -991 -319
rect -933 -1219 -843 -319
rect -785 -1219 -695 -319
rect -637 -1219 -547 -319
rect -489 -1219 -399 -319
rect -341 -1219 -251 -319
rect -193 -1219 -103 -319
rect -45 -1219 45 -319
rect 103 -1219 193 -319
rect 251 -1219 341 -319
rect 399 -1219 489 -319
rect 547 -1219 637 -319
rect 695 -1219 785 -319
rect 843 -1219 933 -319
rect 991 -1219 1081 -319
rect 1139 -1219 1229 -319
rect 1287 -1219 1377 -319
rect 1435 -1219 1525 -319
rect 1583 -1219 1673 -319
rect 1731 -1219 1821 -319
<< pdiff >>
rect -1879 935 -1821 947
rect -1879 59 -1867 935
rect -1833 59 -1821 935
rect -1879 47 -1821 59
rect -1731 935 -1673 947
rect -1731 59 -1719 935
rect -1685 59 -1673 935
rect -1731 47 -1673 59
rect -1583 935 -1525 947
rect -1583 59 -1571 935
rect -1537 59 -1525 935
rect -1583 47 -1525 59
rect -1435 935 -1377 947
rect -1435 59 -1423 935
rect -1389 59 -1377 935
rect -1435 47 -1377 59
rect -1287 935 -1229 947
rect -1287 59 -1275 935
rect -1241 59 -1229 935
rect -1287 47 -1229 59
rect -1139 935 -1081 947
rect -1139 59 -1127 935
rect -1093 59 -1081 935
rect -1139 47 -1081 59
rect -991 935 -933 947
rect -991 59 -979 935
rect -945 59 -933 935
rect -991 47 -933 59
rect -843 935 -785 947
rect -843 59 -831 935
rect -797 59 -785 935
rect -843 47 -785 59
rect -695 935 -637 947
rect -695 59 -683 935
rect -649 59 -637 935
rect -695 47 -637 59
rect -547 935 -489 947
rect -547 59 -535 935
rect -501 59 -489 935
rect -547 47 -489 59
rect -399 935 -341 947
rect -399 59 -387 935
rect -353 59 -341 935
rect -399 47 -341 59
rect -251 935 -193 947
rect -251 59 -239 935
rect -205 59 -193 935
rect -251 47 -193 59
rect -103 935 -45 947
rect -103 59 -91 935
rect -57 59 -45 935
rect -103 47 -45 59
rect 45 935 103 947
rect 45 59 57 935
rect 91 59 103 935
rect 45 47 103 59
rect 193 935 251 947
rect 193 59 205 935
rect 239 59 251 935
rect 193 47 251 59
rect 341 935 399 947
rect 341 59 353 935
rect 387 59 399 935
rect 341 47 399 59
rect 489 935 547 947
rect 489 59 501 935
rect 535 59 547 935
rect 489 47 547 59
rect 637 935 695 947
rect 637 59 649 935
rect 683 59 695 935
rect 637 47 695 59
rect 785 935 843 947
rect 785 59 797 935
rect 831 59 843 935
rect 785 47 843 59
rect 933 935 991 947
rect 933 59 945 935
rect 979 59 991 935
rect 933 47 991 59
rect 1081 935 1139 947
rect 1081 59 1093 935
rect 1127 59 1139 935
rect 1081 47 1139 59
rect 1229 935 1287 947
rect 1229 59 1241 935
rect 1275 59 1287 935
rect 1229 47 1287 59
rect 1377 935 1435 947
rect 1377 59 1389 935
rect 1423 59 1435 935
rect 1377 47 1435 59
rect 1525 935 1583 947
rect 1525 59 1537 935
rect 1571 59 1583 935
rect 1525 47 1583 59
rect 1673 935 1731 947
rect 1673 59 1685 935
rect 1719 59 1731 935
rect 1673 47 1731 59
rect 1821 935 1879 947
rect 1821 59 1833 935
rect 1867 59 1879 935
rect 1821 47 1879 59
rect -1879 -331 -1821 -319
rect -1879 -1207 -1867 -331
rect -1833 -1207 -1821 -331
rect -1879 -1219 -1821 -1207
rect -1731 -331 -1673 -319
rect -1731 -1207 -1719 -331
rect -1685 -1207 -1673 -331
rect -1731 -1219 -1673 -1207
rect -1583 -331 -1525 -319
rect -1583 -1207 -1571 -331
rect -1537 -1207 -1525 -331
rect -1583 -1219 -1525 -1207
rect -1435 -331 -1377 -319
rect -1435 -1207 -1423 -331
rect -1389 -1207 -1377 -331
rect -1435 -1219 -1377 -1207
rect -1287 -331 -1229 -319
rect -1287 -1207 -1275 -331
rect -1241 -1207 -1229 -331
rect -1287 -1219 -1229 -1207
rect -1139 -331 -1081 -319
rect -1139 -1207 -1127 -331
rect -1093 -1207 -1081 -331
rect -1139 -1219 -1081 -1207
rect -991 -331 -933 -319
rect -991 -1207 -979 -331
rect -945 -1207 -933 -331
rect -991 -1219 -933 -1207
rect -843 -331 -785 -319
rect -843 -1207 -831 -331
rect -797 -1207 -785 -331
rect -843 -1219 -785 -1207
rect -695 -331 -637 -319
rect -695 -1207 -683 -331
rect -649 -1207 -637 -331
rect -695 -1219 -637 -1207
rect -547 -331 -489 -319
rect -547 -1207 -535 -331
rect -501 -1207 -489 -331
rect -547 -1219 -489 -1207
rect -399 -331 -341 -319
rect -399 -1207 -387 -331
rect -353 -1207 -341 -331
rect -399 -1219 -341 -1207
rect -251 -331 -193 -319
rect -251 -1207 -239 -331
rect -205 -1207 -193 -331
rect -251 -1219 -193 -1207
rect -103 -331 -45 -319
rect -103 -1207 -91 -331
rect -57 -1207 -45 -331
rect -103 -1219 -45 -1207
rect 45 -331 103 -319
rect 45 -1207 57 -331
rect 91 -1207 103 -331
rect 45 -1219 103 -1207
rect 193 -331 251 -319
rect 193 -1207 205 -331
rect 239 -1207 251 -331
rect 193 -1219 251 -1207
rect 341 -331 399 -319
rect 341 -1207 353 -331
rect 387 -1207 399 -331
rect 341 -1219 399 -1207
rect 489 -331 547 -319
rect 489 -1207 501 -331
rect 535 -1207 547 -331
rect 489 -1219 547 -1207
rect 637 -331 695 -319
rect 637 -1207 649 -331
rect 683 -1207 695 -331
rect 637 -1219 695 -1207
rect 785 -331 843 -319
rect 785 -1207 797 -331
rect 831 -1207 843 -331
rect 785 -1219 843 -1207
rect 933 -331 991 -319
rect 933 -1207 945 -331
rect 979 -1207 991 -331
rect 933 -1219 991 -1207
rect 1081 -331 1139 -319
rect 1081 -1207 1093 -331
rect 1127 -1207 1139 -331
rect 1081 -1219 1139 -1207
rect 1229 -331 1287 -319
rect 1229 -1207 1241 -331
rect 1275 -1207 1287 -331
rect 1229 -1219 1287 -1207
rect 1377 -331 1435 -319
rect 1377 -1207 1389 -331
rect 1423 -1207 1435 -331
rect 1377 -1219 1435 -1207
rect 1525 -331 1583 -319
rect 1525 -1207 1537 -331
rect 1571 -1207 1583 -331
rect 1525 -1219 1583 -1207
rect 1673 -331 1731 -319
rect 1673 -1207 1685 -331
rect 1719 -1207 1731 -331
rect 1673 -1219 1731 -1207
rect 1821 -331 1879 -319
rect 1821 -1207 1833 -331
rect 1867 -1207 1879 -331
rect 1821 -1219 1879 -1207
<< pdiffc >>
rect -1867 59 -1833 935
rect -1719 59 -1685 935
rect -1571 59 -1537 935
rect -1423 59 -1389 935
rect -1275 59 -1241 935
rect -1127 59 -1093 935
rect -979 59 -945 935
rect -831 59 -797 935
rect -683 59 -649 935
rect -535 59 -501 935
rect -387 59 -353 935
rect -239 59 -205 935
rect -91 59 -57 935
rect 57 59 91 935
rect 205 59 239 935
rect 353 59 387 935
rect 501 59 535 935
rect 649 59 683 935
rect 797 59 831 935
rect 945 59 979 935
rect 1093 59 1127 935
rect 1241 59 1275 935
rect 1389 59 1423 935
rect 1537 59 1571 935
rect 1685 59 1719 935
rect 1833 59 1867 935
rect -1867 -1207 -1833 -331
rect -1719 -1207 -1685 -331
rect -1571 -1207 -1537 -331
rect -1423 -1207 -1389 -331
rect -1275 -1207 -1241 -331
rect -1127 -1207 -1093 -331
rect -979 -1207 -945 -331
rect -831 -1207 -797 -331
rect -683 -1207 -649 -331
rect -535 -1207 -501 -331
rect -387 -1207 -353 -331
rect -239 -1207 -205 -331
rect -91 -1207 -57 -331
rect 57 -1207 91 -331
rect 205 -1207 239 -331
rect 353 -1207 387 -331
rect 501 -1207 535 -331
rect 649 -1207 683 -331
rect 797 -1207 831 -331
rect 945 -1207 979 -331
rect 1093 -1207 1127 -331
rect 1241 -1207 1275 -331
rect 1389 -1207 1423 -331
rect 1537 -1207 1571 -331
rect 1685 -1207 1719 -331
rect 1833 -1207 1867 -331
<< nsubdiff >>
rect -1947 1126 -1885 1160
rect 1885 1126 1947 1160
rect -1947 1025 -1885 1059
rect 1885 1025 1947 1059
<< nsubdiffcont >>
rect -1885 1126 1885 1160
rect -1885 1025 1885 1059
<< poly >>
rect -2017 964 2017 1005
rect -1821 947 -1731 964
rect -1673 947 -1583 964
rect -1525 947 -1435 964
rect -1377 947 -1287 964
rect -1229 947 -1139 964
rect -1081 947 -991 964
rect -933 947 -843 964
rect -785 947 -695 964
rect -637 947 -547 964
rect -489 947 -399 964
rect -341 947 -251 964
rect -193 947 -103 964
rect -45 947 45 964
rect 103 947 193 964
rect 251 947 341 964
rect 399 947 489 964
rect 547 947 637 964
rect 695 947 785 964
rect 843 947 933 964
rect 991 947 1081 964
rect 1139 947 1229 964
rect 1287 947 1377 964
rect 1435 947 1525 964
rect 1583 947 1673 964
rect 1731 947 1821 964
rect -1821 24 -1731 47
rect -1673 24 -1583 47
rect -1525 24 -1435 47
rect -1377 24 -1287 47
rect -1229 24 -1139 47
rect -1081 24 -991 47
rect -933 24 -843 47
rect -785 24 -695 47
rect -637 24 -547 47
rect -489 24 -399 47
rect -341 24 -251 47
rect -193 24 -103 47
rect -45 24 45 47
rect 103 24 193 47
rect 251 24 341 47
rect 399 24 489 47
rect 547 24 637 47
rect 695 24 785 47
rect 843 24 933 47
rect 991 24 1081 47
rect 1139 24 1229 47
rect 1287 24 1377 47
rect 1435 24 1525 47
rect 1583 24 1673 47
rect 1731 24 1821 47
rect -2017 -10 2017 24
rect -2017 -44 -1902 -10
rect -1778 -44 -1610 -10
rect -1486 -44 -1303 -10
rect -1179 -44 -1027 -10
rect -903 -44 -720 -10
rect -596 -44 -413 -10
rect -289 -44 -137 -10
rect -13 -44 170 -10
rect 294 -44 447 -10
rect 571 -44 767 -10
rect 891 -44 1040 -10
rect 1164 -44 1342 -10
rect 1466 -44 1645 -10
rect 1769 -44 2017 -10
rect -2017 -61 2017 -44
rect -2017 -230 2017 -211
rect -2017 -264 -1903 -230
rect -1779 -264 -1616 -230
rect -1492 -264 -1312 -230
rect -1188 -264 -1007 -230
rect -883 -264 -738 -230
rect -614 -264 -433 -230
rect -309 -264 -128 -230
rect -4 -264 176 -230
rect 300 -264 463 -230
rect 587 -264 768 -230
rect 892 -264 1046 -230
rect 1170 -264 1351 -230
rect 1475 -264 1656 -230
rect 1780 -264 2017 -230
rect -2017 -295 2017 -264
rect -1821 -319 -1731 -295
rect -1673 -319 -1583 -295
rect -1525 -319 -1435 -295
rect -1377 -319 -1287 -295
rect -1229 -319 -1139 -295
rect -1081 -319 -991 -295
rect -933 -319 -843 -295
rect -785 -319 -695 -295
rect -637 -319 -547 -295
rect -489 -319 -399 -295
rect -341 -319 -251 -295
rect -193 -319 -103 -295
rect -45 -319 45 -295
rect 103 -319 193 -295
rect 251 -319 341 -295
rect 399 -319 489 -295
rect 547 -319 637 -295
rect 695 -319 785 -295
rect 843 -319 933 -295
rect 991 -319 1081 -295
rect 1139 -319 1229 -295
rect 1287 -319 1377 -295
rect 1435 -319 1525 -295
rect 1583 -319 1673 -295
rect 1731 -319 1821 -295
rect -1821 -1241 -1731 -1219
rect -1673 -1241 -1583 -1219
rect -1525 -1241 -1435 -1219
rect -1377 -1241 -1287 -1219
rect -1229 -1241 -1139 -1219
rect -1081 -1241 -991 -1219
rect -933 -1241 -843 -1219
rect -785 -1241 -695 -1219
rect -637 -1241 -547 -1219
rect -489 -1241 -399 -1219
rect -341 -1241 -251 -1219
rect -193 -1241 -103 -1219
rect -45 -1241 45 -1219
rect 103 -1241 193 -1219
rect 251 -1241 341 -1219
rect 399 -1241 489 -1219
rect 547 -1241 637 -1219
rect 695 -1241 785 -1219
rect 843 -1241 933 -1219
rect 991 -1241 1081 -1219
rect 1139 -1241 1229 -1219
rect 1287 -1241 1377 -1219
rect 1435 -1241 1525 -1219
rect 1583 -1241 1673 -1219
rect 1731 -1241 1821 -1219
rect -2017 -1317 2017 -1241
<< polycont >>
rect -1902 -44 -1778 -10
rect -1610 -44 -1486 -10
rect -1303 -44 -1179 -10
rect -1027 -44 -903 -10
rect -720 -44 -596 -10
rect -413 -44 -289 -10
rect -137 -44 -13 -10
rect 170 -44 294 -10
rect 447 -44 571 -10
rect 767 -44 891 -10
rect 1040 -44 1164 -10
rect 1342 -44 1466 -10
rect 1645 -44 1769 -10
rect -1903 -264 -1779 -230
rect -1616 -264 -1492 -230
rect -1312 -264 -1188 -230
rect -1007 -264 -883 -230
rect -738 -264 -614 -230
rect -433 -264 -309 -230
rect -128 -264 -4 -230
rect 176 -264 300 -230
rect 463 -264 587 -230
rect 768 -264 892 -230
rect 1046 -264 1170 -230
rect 1351 -264 1475 -230
rect 1656 -264 1780 -230
<< locali >>
rect -1947 1126 -1885 1160
rect 1885 1126 1947 1160
rect -1947 1025 -1885 1059
rect 1885 1025 1947 1059
rect -1867 935 -1833 951
rect -1867 43 -1833 59
rect -1719 935 -1685 951
rect -1719 43 -1685 59
rect -1571 935 -1537 951
rect -1571 43 -1537 59
rect -1423 935 -1389 951
rect -1423 43 -1389 59
rect -1275 935 -1241 951
rect -1275 43 -1241 59
rect -1127 935 -1093 951
rect -1127 43 -1093 59
rect -979 935 -945 951
rect -979 43 -945 59
rect -831 935 -797 951
rect -831 43 -797 59
rect -683 935 -649 951
rect -683 43 -649 59
rect -535 935 -501 951
rect -535 43 -501 59
rect -387 935 -353 951
rect -387 43 -353 59
rect -239 935 -205 951
rect -239 43 -205 59
rect -91 935 -57 951
rect -91 43 -57 59
rect 57 935 91 951
rect 57 43 91 59
rect 205 935 239 951
rect 205 43 239 59
rect 353 935 387 951
rect 353 43 387 59
rect 501 935 535 951
rect 501 43 535 59
rect 649 935 683 951
rect 649 43 683 59
rect 797 935 831 951
rect 797 43 831 59
rect 945 935 979 951
rect 945 43 979 59
rect 1093 935 1127 951
rect 1093 43 1127 59
rect 1241 935 1275 951
rect 1241 43 1275 59
rect 1389 935 1423 951
rect 1389 43 1423 59
rect 1537 935 1571 951
rect 1537 43 1571 59
rect 1685 935 1719 951
rect 1685 43 1719 59
rect 1833 935 1867 951
rect 1833 43 1867 59
rect -1918 -10 -1761 7
rect -1918 -44 -1902 -10
rect -1778 -44 -1761 -10
rect -1918 -61 -1761 -44
rect -1626 -10 -1469 7
rect -1626 -44 -1610 -10
rect -1486 -44 -1469 -10
rect -1626 -61 -1469 -44
rect -1319 -10 -1162 7
rect -1319 -44 -1303 -10
rect -1179 -44 -1162 -10
rect -1319 -61 -1162 -44
rect -1043 -10 -886 7
rect -1043 -44 -1027 -10
rect -903 -44 -886 -10
rect -1043 -61 -886 -44
rect -736 -10 -579 7
rect -736 -44 -720 -10
rect -596 -44 -579 -10
rect -736 -61 -579 -44
rect -429 -10 -272 7
rect -429 -44 -413 -10
rect -289 -44 -272 -10
rect -429 -61 -272 -44
rect -153 -10 4 7
rect -153 -44 -137 -10
rect -13 -44 4 -10
rect -153 -61 4 -44
rect 154 -10 311 7
rect 154 -44 170 -10
rect 294 -44 311 -10
rect 154 -61 311 -44
rect 431 -10 588 7
rect 431 -44 447 -10
rect 571 -44 588 -10
rect 431 -61 588 -44
rect 751 -10 908 7
rect 751 -44 767 -10
rect 891 -44 908 -10
rect 751 -61 908 -44
rect 1024 -10 1181 7
rect 1024 -44 1040 -10
rect 1164 -44 1181 -10
rect 1024 -61 1181 -44
rect 1326 -10 1483 7
rect 1326 -44 1342 -10
rect 1466 -44 1483 -10
rect 1326 -61 1483 -44
rect 1629 -10 1786 7
rect 1629 -44 1645 -10
rect 1769 -44 1786 -10
rect 1629 -61 1786 -44
rect -1919 -230 -1763 -213
rect -1919 -264 -1903 -230
rect -1779 -264 -1763 -230
rect -1919 -281 -1763 -264
rect -1632 -230 -1476 -213
rect -1632 -264 -1616 -230
rect -1492 -264 -1476 -230
rect -1632 -281 -1476 -264
rect -1328 -230 -1172 -213
rect -1328 -264 -1312 -230
rect -1188 -264 -1172 -230
rect -1328 -281 -1172 -264
rect -1023 -230 -867 -213
rect -1023 -264 -1007 -230
rect -883 -264 -867 -230
rect -1023 -281 -867 -264
rect -754 -230 -598 -213
rect -754 -264 -738 -230
rect -614 -264 -598 -230
rect -754 -281 -598 -264
rect -449 -230 -293 -213
rect -449 -264 -433 -230
rect -309 -264 -293 -230
rect -449 -281 -293 -264
rect -144 -230 12 -213
rect -144 -264 -128 -230
rect -4 -264 12 -230
rect -144 -281 12 -264
rect 160 -230 316 -213
rect 160 -264 176 -230
rect 300 -264 316 -230
rect 160 -281 316 -264
rect 447 -230 603 -213
rect 447 -264 463 -230
rect 587 -264 603 -230
rect 447 -281 603 -264
rect 752 -230 908 -213
rect 752 -264 768 -230
rect 892 -264 908 -230
rect 752 -281 908 -264
rect 1030 -230 1186 -213
rect 1030 -264 1046 -230
rect 1170 -264 1186 -230
rect 1030 -281 1186 -264
rect 1335 -230 1491 -213
rect 1335 -264 1351 -230
rect 1475 -264 1491 -230
rect 1335 -281 1491 -264
rect 1640 -230 1796 -213
rect 1640 -264 1656 -230
rect 1780 -264 1796 -230
rect 1640 -281 1796 -264
rect -1867 -331 -1833 -315
rect -1867 -1223 -1833 -1207
rect -1719 -331 -1685 -315
rect -1719 -1223 -1685 -1207
rect -1571 -331 -1537 -315
rect -1571 -1223 -1537 -1207
rect -1423 -331 -1389 -315
rect -1423 -1223 -1389 -1207
rect -1275 -331 -1241 -315
rect -1275 -1223 -1241 -1207
rect -1127 -331 -1093 -315
rect -1127 -1223 -1093 -1207
rect -979 -331 -945 -315
rect -979 -1223 -945 -1207
rect -831 -331 -797 -315
rect -831 -1223 -797 -1207
rect -683 -331 -649 -315
rect -683 -1223 -649 -1207
rect -535 -331 -501 -315
rect -535 -1223 -501 -1207
rect -387 -331 -353 -315
rect -387 -1223 -353 -1207
rect -239 -331 -205 -315
rect -239 -1223 -205 -1207
rect -91 -331 -57 -315
rect -91 -1223 -57 -1207
rect 57 -331 91 -315
rect 57 -1223 91 -1207
rect 205 -331 239 -315
rect 205 -1223 239 -1207
rect 353 -331 387 -315
rect 353 -1223 387 -1207
rect 501 -331 535 -315
rect 501 -1223 535 -1207
rect 649 -331 683 -315
rect 649 -1223 683 -1207
rect 797 -331 831 -315
rect 797 -1223 831 -1207
rect 945 -331 979 -315
rect 945 -1223 979 -1207
rect 1093 -331 1127 -315
rect 1093 -1223 1127 -1207
rect 1241 -331 1275 -315
rect 1241 -1223 1275 -1207
rect 1389 -331 1423 -315
rect 1389 -1223 1423 -1207
rect 1537 -331 1571 -315
rect 1537 -1223 1571 -1207
rect 1685 -331 1719 -315
rect 1685 -1223 1719 -1207
rect 1833 -331 1867 -315
rect 1833 -1223 1867 -1207
<< viali >>
rect -1885 1126 1885 1160
rect -1885 1025 1885 1059
rect -1867 59 -1833 935
rect -1719 59 -1685 935
rect -1571 59 -1537 935
rect -1423 59 -1389 935
rect -1275 59 -1241 935
rect -1127 59 -1093 935
rect -979 59 -945 935
rect -831 59 -797 935
rect -683 59 -649 935
rect -535 59 -501 935
rect -387 59 -353 935
rect -239 59 -205 935
rect -91 59 -57 935
rect 57 59 91 935
rect 205 59 239 935
rect 353 59 387 935
rect 501 59 535 935
rect 649 59 683 935
rect 797 59 831 935
rect 945 59 979 935
rect 1093 59 1127 935
rect 1241 59 1275 935
rect 1389 59 1423 935
rect 1537 59 1571 935
rect 1685 59 1719 935
rect 1833 59 1867 935
rect -1902 -44 -1778 -10
rect -1610 -44 -1486 -10
rect -1303 -44 -1179 -10
rect -1027 -44 -903 -10
rect -720 -44 -596 -10
rect -413 -44 -289 -10
rect -137 -44 -13 -10
rect 170 -44 294 -10
rect 447 -44 571 -10
rect 767 -44 891 -10
rect 1040 -44 1164 -10
rect 1342 -44 1466 -10
rect 1645 -44 1769 -10
rect -1903 -264 -1779 -230
rect -1616 -264 -1492 -230
rect -1312 -264 -1188 -230
rect -1007 -264 -883 -230
rect -738 -264 -614 -230
rect -433 -264 -309 -230
rect -128 -264 -4 -230
rect 176 -264 300 -230
rect 463 -264 587 -230
rect 768 -264 892 -230
rect 1046 -264 1170 -230
rect 1351 -264 1475 -230
rect 1656 -264 1780 -230
rect -1867 -1207 -1833 -331
rect -1719 -1207 -1685 -331
rect -1571 -1207 -1537 -331
rect -1423 -1207 -1389 -331
rect -1275 -1207 -1241 -331
rect -1127 -1207 -1093 -331
rect -979 -1207 -945 -331
rect -831 -1207 -797 -331
rect -683 -1207 -649 -331
rect -535 -1207 -501 -331
rect -387 -1207 -353 -331
rect -239 -1207 -205 -331
rect -91 -1207 -57 -331
rect 57 -1207 91 -331
rect 205 -1207 239 -331
rect 353 -1207 387 -331
rect 501 -1207 535 -331
rect 649 -1207 683 -331
rect 797 -1207 831 -331
rect 945 -1207 979 -331
rect 1093 -1207 1127 -331
rect 1241 -1207 1275 -331
rect 1389 -1207 1423 -331
rect 1537 -1207 1571 -331
rect 1685 -1207 1719 -331
rect 1833 -1207 1867 -331
<< metal1 >>
rect -2017 1160 2017 1167
rect -2017 1126 -1885 1160
rect 1885 1126 2017 1160
rect -2017 1059 2017 1126
rect -2017 1025 -1885 1059
rect 1885 1025 2017 1059
rect -2017 1018 2017 1025
rect -1873 935 -1827 1018
rect -1873 59 -1867 935
rect -1833 59 -1827 935
rect -1873 46 -1827 59
rect -1725 935 -1679 947
rect -1725 59 -1719 935
rect -1685 59 -1679 935
rect -1923 -55 -1913 0
rect -1773 -55 -1763 0
rect -1725 -99 -1679 59
rect -1577 935 -1531 1018
rect -1577 59 -1571 935
rect -1537 59 -1531 935
rect -1577 47 -1531 59
rect -1429 935 -1383 947
rect -1429 59 -1423 935
rect -1389 59 -1383 935
rect -1631 -55 -1621 0
rect -1481 -55 -1471 0
rect -1429 -99 -1383 59
rect -1281 935 -1235 1018
rect -986 947 -940 1018
rect -1281 59 -1275 935
rect -1241 59 -1235 935
rect -1281 46 -1235 59
rect -1133 935 -1087 947
rect -1133 59 -1127 935
rect -1093 59 -1087 935
rect -1324 -55 -1314 0
rect -1174 -55 -1164 0
rect -1133 -99 -1087 59
rect -986 935 -939 947
rect -986 59 -979 935
rect -945 59 -939 935
rect -986 47 -939 59
rect -837 935 -791 947
rect -837 59 -831 935
rect -797 59 -791 935
rect -986 46 -940 47
rect -1048 -55 -1038 0
rect -898 -55 -888 0
rect -837 -99 -791 59
rect -689 935 -643 1018
rect -689 59 -683 935
rect -649 59 -643 935
rect -689 46 -643 59
rect -541 935 -495 947
rect -541 59 -535 935
rect -501 59 -495 935
rect -741 -55 -731 0
rect -591 -55 -581 0
rect -541 -99 -495 59
rect -393 935 -347 1018
rect -393 59 -387 935
rect -353 59 -347 935
rect -393 47 -347 59
rect -245 935 -199 947
rect -245 59 -239 935
rect -205 59 -199 935
rect -434 -55 -424 0
rect -284 -55 -274 0
rect -245 -99 -199 59
rect -97 935 -51 1018
rect -97 59 -91 935
rect -57 59 -51 935
rect -97 47 -51 59
rect 51 935 97 947
rect 51 59 57 935
rect 91 59 97 935
rect -158 -55 -148 0
rect -8 -55 2 0
rect 51 -99 97 59
rect 199 935 245 1018
rect 199 59 205 935
rect 239 59 245 935
rect 199 47 245 59
rect 347 935 393 947
rect 347 59 353 935
rect 387 59 393 935
rect 149 -55 159 0
rect 299 -55 309 0
rect 347 -99 393 59
rect 495 935 541 1018
rect 495 59 501 935
rect 535 59 541 935
rect 495 46 541 59
rect 643 935 689 947
rect 643 59 649 935
rect 683 59 689 935
rect 426 -55 436 0
rect 576 -55 586 0
rect 643 -99 689 59
rect 791 935 837 1018
rect 791 59 797 935
rect 831 59 837 935
rect 791 46 837 59
rect 939 935 985 947
rect 939 59 945 935
rect 979 59 985 935
rect 746 -55 756 0
rect 896 -55 906 0
rect 939 -99 985 59
rect 1087 935 1133 1018
rect 1087 59 1093 935
rect 1127 59 1133 935
rect 1087 46 1133 59
rect 1235 935 1281 947
rect 1235 59 1241 935
rect 1275 59 1281 935
rect 1019 -55 1029 0
rect 1169 -55 1179 0
rect 1235 -99 1281 59
rect 1383 935 1429 1018
rect 1383 59 1389 935
rect 1423 59 1429 935
rect 1383 46 1429 59
rect 1531 935 1577 947
rect 1531 59 1537 935
rect 1571 59 1577 935
rect 1321 -55 1331 0
rect 1471 -55 1481 0
rect 1531 -99 1577 59
rect 1679 935 1725 1018
rect 1679 59 1685 935
rect 1719 59 1725 935
rect 1679 47 1725 59
rect 1827 935 1873 947
rect 1827 59 1833 935
rect 1867 59 1873 935
rect 1624 -55 1634 0
rect 1774 -55 1784 0
rect 1827 -99 1873 59
rect -1725 -170 1873 -99
rect -1919 -271 -1909 -219
rect -1777 -271 -1767 -219
rect -1873 -331 -1827 -319
rect -1873 -1207 -1867 -331
rect -1833 -1207 -1827 -331
rect -1873 -1315 -1827 -1207
rect -1725 -331 -1679 -170
rect -1632 -271 -1622 -219
rect -1490 -271 -1480 -219
rect -1725 -1207 -1719 -331
rect -1685 -1207 -1679 -331
rect -1725 -1219 -1679 -1207
rect -1577 -331 -1531 -319
rect -1577 -1207 -1571 -331
rect -1537 -1207 -1531 -331
rect -1577 -1315 -1531 -1207
rect -1429 -331 -1383 -170
rect -1328 -271 -1318 -219
rect -1186 -271 -1176 -219
rect -1429 -1207 -1423 -331
rect -1389 -1207 -1383 -331
rect -1429 -1219 -1383 -1207
rect -1281 -331 -1235 -319
rect -1281 -1207 -1275 -331
rect -1241 -1207 -1235 -331
rect -1281 -1315 -1235 -1207
rect -1133 -331 -1087 -170
rect -1023 -271 -1013 -219
rect -881 -271 -871 -219
rect -1133 -1207 -1127 -331
rect -1093 -1207 -1087 -331
rect -1133 -1219 -1087 -1207
rect -985 -331 -939 -319
rect -985 -1207 -979 -331
rect -945 -1207 -939 -331
rect -985 -1315 -939 -1207
rect -837 -331 -791 -170
rect -754 -271 -744 -219
rect -612 -271 -602 -219
rect -837 -1207 -831 -331
rect -797 -1207 -791 -331
rect -837 -1219 -791 -1207
rect -689 -331 -643 -319
rect -689 -1207 -683 -331
rect -649 -1207 -643 -331
rect -689 -1315 -643 -1207
rect -541 -331 -495 -170
rect -449 -271 -439 -219
rect -307 -271 -297 -219
rect -541 -1207 -535 -331
rect -501 -1207 -495 -331
rect -541 -1219 -495 -1207
rect -393 -331 -347 -319
rect -393 -1207 -387 -331
rect -353 -1207 -347 -331
rect -393 -1315 -347 -1207
rect -245 -331 -199 -170
rect -144 -271 -134 -219
rect -2 -271 8 -219
rect -245 -1207 -239 -331
rect -205 -1207 -199 -331
rect -245 -1219 -199 -1207
rect -97 -331 -51 -319
rect -97 -1207 -91 -331
rect -57 -1207 -51 -331
rect -97 -1315 -51 -1207
rect 51 -331 97 -170
rect 160 -271 170 -219
rect 302 -271 312 -219
rect 51 -1207 57 -331
rect 91 -1207 97 -331
rect 51 -1219 97 -1207
rect 199 -331 245 -319
rect 199 -1207 205 -331
rect 239 -1207 245 -331
rect 199 -1315 245 -1207
rect 347 -331 393 -170
rect 447 -271 457 -219
rect 589 -271 599 -219
rect 347 -1207 353 -331
rect 387 -1207 393 -331
rect 347 -1219 393 -1207
rect 495 -331 541 -319
rect 495 -1207 501 -331
rect 535 -1207 541 -331
rect 495 -1315 541 -1207
rect 643 -331 689 -170
rect 752 -271 762 -219
rect 894 -271 904 -219
rect 643 -1207 649 -331
rect 683 -1207 689 -331
rect 643 -1219 689 -1207
rect 791 -331 837 -319
rect 791 -1207 797 -331
rect 831 -1207 837 -331
rect 791 -1315 837 -1207
rect 939 -331 985 -170
rect 1030 -271 1040 -219
rect 1172 -271 1182 -219
rect 939 -1207 945 -331
rect 979 -1207 985 -331
rect 939 -1219 985 -1207
rect 1087 -331 1133 -319
rect 1087 -1207 1093 -331
rect 1127 -1207 1133 -331
rect 1087 -1315 1133 -1207
rect 1235 -331 1281 -170
rect 1335 -271 1345 -219
rect 1477 -271 1487 -219
rect 1235 -1207 1241 -331
rect 1275 -1207 1281 -331
rect 1235 -1219 1281 -1207
rect 1383 -331 1429 -319
rect 1383 -1207 1389 -331
rect 1423 -1207 1429 -331
rect 1383 -1315 1429 -1207
rect 1531 -331 1577 -170
rect 1640 -271 1650 -219
rect 1782 -271 1792 -219
rect 1531 -1207 1537 -331
rect 1571 -1207 1577 -331
rect 1531 -1219 1577 -1207
rect 1679 -331 1725 -319
rect 1679 -1207 1685 -331
rect 1719 -1207 1725 -331
rect 1679 -1315 1725 -1207
rect 1827 -331 1873 -170
rect 1827 -1207 1833 -331
rect 1867 -1207 1873 -331
rect 1827 -1219 1873 -1207
rect -1950 -1454 1949 -1315
<< via1 >>
rect -1913 -10 -1773 0
rect -1913 -44 -1902 -10
rect -1902 -44 -1778 -10
rect -1778 -44 -1773 -10
rect -1913 -55 -1773 -44
rect -1621 -10 -1481 0
rect -1621 -44 -1610 -10
rect -1610 -44 -1486 -10
rect -1486 -44 -1481 -10
rect -1621 -55 -1481 -44
rect -1314 -10 -1174 0
rect -1314 -44 -1303 -10
rect -1303 -44 -1179 -10
rect -1179 -44 -1174 -10
rect -1314 -55 -1174 -44
rect -1038 -10 -898 0
rect -1038 -44 -1027 -10
rect -1027 -44 -903 -10
rect -903 -44 -898 -10
rect -1038 -55 -898 -44
rect -731 -10 -591 0
rect -731 -44 -720 -10
rect -720 -44 -596 -10
rect -596 -44 -591 -10
rect -731 -55 -591 -44
rect -424 -10 -284 0
rect -424 -44 -413 -10
rect -413 -44 -289 -10
rect -289 -44 -284 -10
rect -424 -55 -284 -44
rect -148 -10 -8 0
rect -148 -44 -137 -10
rect -137 -44 -13 -10
rect -13 -44 -8 -10
rect -148 -55 -8 -44
rect 159 -10 299 0
rect 159 -44 170 -10
rect 170 -44 294 -10
rect 294 -44 299 -10
rect 159 -55 299 -44
rect 436 -10 576 0
rect 436 -44 447 -10
rect 447 -44 571 -10
rect 571 -44 576 -10
rect 436 -55 576 -44
rect 756 -10 896 0
rect 756 -44 767 -10
rect 767 -44 891 -10
rect 891 -44 896 -10
rect 756 -55 896 -44
rect 1029 -10 1169 0
rect 1029 -44 1040 -10
rect 1040 -44 1164 -10
rect 1164 -44 1169 -10
rect 1029 -55 1169 -44
rect 1331 -10 1471 0
rect 1331 -44 1342 -10
rect 1342 -44 1466 -10
rect 1466 -44 1471 -10
rect 1331 -55 1471 -44
rect 1634 -10 1774 0
rect 1634 -44 1645 -10
rect 1645 -44 1769 -10
rect 1769 -44 1774 -10
rect 1634 -55 1774 -44
rect -1909 -230 -1777 -219
rect -1909 -264 -1903 -230
rect -1903 -264 -1779 -230
rect -1779 -264 -1777 -230
rect -1909 -271 -1777 -264
rect -1622 -230 -1490 -219
rect -1622 -264 -1616 -230
rect -1616 -264 -1492 -230
rect -1492 -264 -1490 -230
rect -1622 -271 -1490 -264
rect -1318 -230 -1186 -219
rect -1318 -264 -1312 -230
rect -1312 -264 -1188 -230
rect -1188 -264 -1186 -230
rect -1318 -271 -1186 -264
rect -1013 -230 -881 -219
rect -1013 -264 -1007 -230
rect -1007 -264 -883 -230
rect -883 -264 -881 -230
rect -1013 -271 -881 -264
rect -744 -230 -612 -219
rect -744 -264 -738 -230
rect -738 -264 -614 -230
rect -614 -264 -612 -230
rect -744 -271 -612 -264
rect -439 -230 -307 -219
rect -439 -264 -433 -230
rect -433 -264 -309 -230
rect -309 -264 -307 -230
rect -439 -271 -307 -264
rect -134 -230 -2 -219
rect -134 -264 -128 -230
rect -128 -264 -4 -230
rect -4 -264 -2 -230
rect -134 -271 -2 -264
rect 170 -230 302 -219
rect 170 -264 176 -230
rect 176 -264 300 -230
rect 300 -264 302 -230
rect 170 -271 302 -264
rect 457 -230 589 -219
rect 457 -264 463 -230
rect 463 -264 587 -230
rect 587 -264 589 -230
rect 457 -271 589 -264
rect 762 -230 894 -219
rect 762 -264 768 -230
rect 768 -264 892 -230
rect 892 -264 894 -230
rect 762 -271 894 -264
rect 1040 -230 1172 -219
rect 1040 -264 1046 -230
rect 1046 -264 1170 -230
rect 1170 -264 1172 -230
rect 1040 -271 1172 -264
rect 1345 -230 1477 -219
rect 1345 -264 1351 -230
rect 1351 -264 1475 -230
rect 1475 -264 1477 -230
rect 1345 -271 1477 -264
rect 1650 -230 1782 -219
rect 1650 -264 1656 -230
rect 1656 -264 1780 -230
rect 1780 -264 1782 -230
rect 1650 -271 1782 -264
<< metal2 >>
rect -2017 0 2017 13
rect -2017 -55 -1913 0
rect -1773 -55 -1621 0
rect -1481 -55 -1314 0
rect -1174 -55 -1038 0
rect -898 -55 -731 0
rect -591 -55 -424 0
rect -284 -55 -148 0
rect -8 -55 159 0
rect 299 -55 436 0
rect 576 -55 756 0
rect 896 -55 1029 0
rect 1169 -55 1331 0
rect 1471 -55 1634 0
rect 1774 -55 2017 0
rect -2017 -57 2017 -55
rect -1913 -65 -1773 -57
rect -1621 -65 -1481 -57
rect -1314 -65 -1174 -57
rect -1038 -65 -898 -57
rect -731 -65 -591 -57
rect -424 -65 -284 -57
rect -148 -65 -8 -57
rect 159 -65 299 -57
rect 436 -65 576 -57
rect 756 -65 896 -57
rect 1029 -65 1169 -57
rect 1331 -65 1471 -57
rect 1634 -65 1774 -57
rect -1909 -215 -1777 -209
rect -1622 -215 -1490 -209
rect -1318 -215 -1186 -209
rect -1013 -215 -881 -209
rect -744 -215 -612 -209
rect -439 -215 -307 -209
rect -134 -215 -2 -209
rect 170 -215 302 -209
rect 457 -215 589 -209
rect 762 -215 894 -209
rect 1040 -215 1172 -209
rect 1345 -215 1477 -209
rect 1650 -215 1782 -209
rect -2017 -219 2017 -215
rect -2017 -271 -1909 -219
rect -1777 -271 -1622 -219
rect -1490 -271 -1318 -219
rect -1186 -271 -1013 -219
rect -881 -271 -744 -219
rect -612 -271 -439 -219
rect -307 -271 -134 -219
rect -2 -271 170 -219
rect 302 -271 457 -219
rect 589 -271 762 -219
rect 894 -271 1040 -219
rect 1172 -271 1345 -219
rect 1477 -271 1650 -219
rect 1782 -271 2017 -219
rect -2017 -285 2017 -271
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -1964 -1042 1964 1042
string parameters w 4.5 l 0.45 m 2 nf 25 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
