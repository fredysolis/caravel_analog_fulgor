* NGSPICE file created from top_pll_v3.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_4ML9WA VSUBS a_429_n486# w_n2457_n634# a_887_n486#
+ a_n29_n486# a_1345_n486# a_n2261_n512# a_1803_n486# a_n487_n486# a_n945_n486# a_n2319_n486#
+ a_n1403_n486# a_2261_n486# a_n1861_n486#
X0 a_2261_n486# a_n2261_n512# a_1803_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X1 a_n945_n486# a_n2261_n512# a_n1403_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X2 a_429_n486# a_n2261_n512# a_n29_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X3 a_1803_n486# a_n2261_n512# a_1345_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X4 a_887_n486# a_n2261_n512# a_429_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X5 a_n487_n486# a_n2261_n512# a_n945_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X6 a_n1403_n486# a_n2261_n512# a_n1861_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X7 a_n1861_n486# a_n2261_n512# a_n2319_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X8 a_n29_n486# a_n2261_n512# a_n487_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X9 a_1345_n486# a_n2261_n512# a_887_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
C0 a_n2319_n486# w_n2457_n634# 0.02fF
C1 a_429_n486# w_n2457_n634# 0.02fF
C2 a_n1403_n486# w_n2457_n634# 0.02fF
C3 w_n2457_n634# a_2261_n486# 0.02fF
C4 w_n2457_n634# a_n1861_n486# 0.02fF
C5 w_n2457_n634# a_n945_n486# 0.02fF
C6 a_1803_n486# w_n2457_n634# 0.02fF
C7 w_n2457_n634# a_n29_n486# 0.02fF
C8 w_n2457_n634# a_n487_n486# 0.02fF
C9 w_n2457_n634# a_1345_n486# 0.02fF
C10 a_887_n486# w_n2457_n634# 0.02fF
C11 a_2261_n486# VSUBS 0.03fF
C12 a_1803_n486# VSUBS 0.03fF
C13 a_1345_n486# VSUBS 0.03fF
C14 a_887_n486# VSUBS 0.03fF
C15 a_429_n486# VSUBS 0.03fF
C16 a_n29_n486# VSUBS 0.03fF
C17 a_n487_n486# VSUBS 0.03fF
C18 a_n945_n486# VSUBS 0.03fF
C19 a_n1403_n486# VSUBS 0.03fF
C20 a_n1861_n486# VSUBS 0.03fF
C21 a_n2319_n486# VSUBS 0.03fF
C22 a_n2261_n512# VSUBS 4.27fF
C23 w_n2457_n634# VSUBS 21.34fF
.ends

.subckt sky130_fd_pr__nfet_01v8_YCGG98 a_n1041_n75# a_n561_n75# a_1167_n75# a_303_n75#
+ a_687_n75# a_n849_n75# a_n369_n75# a_975_n75# a_111_n75# a_495_n75# a_n1137_n75#
+ a_n657_n75# a_n177_n75# a_783_n75# a_n945_n75# a_n465_n75# a_207_n75# a_1071_n75#
+ a_591_n75# a_15_n75# a_n753_n75# w_n1367_n285# a_n273_n75# a_879_n75# a_399_n75#
+ a_n1229_n75# a_n81_n75# a_n1167_n101#
X0 a_207_n75# a_n1167_n101# a_111_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_303_n75# a_n1167_n101# a_207_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_399_n75# a_n1167_n101# a_303_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_495_n75# a_n1167_n101# a_399_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_591_n75# a_n1167_n101# a_495_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_783_n75# a_n1167_n101# a_687_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_687_n75# a_n1167_n101# a_591_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_879_n75# a_n1167_n101# a_783_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_975_n75# a_n1167_n101# a_879_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_n1041_n75# a_n1167_n101# a_n1137_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_n1137_n75# a_n1167_n101# a_n1229_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n561_n75# a_n1167_n101# a_n657_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_1071_n75# a_n1167_n101# a_975_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n945_n75# a_n1167_n101# a_n1041_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n753_n75# a_n1167_n101# a_n849_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n657_n75# a_n1167_n101# a_n753_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n465_n75# a_n1167_n101# a_n561_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n369_n75# a_n1167_n101# a_n465_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_1167_n75# a_n1167_n101# a_1071_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n849_n75# a_n1167_n101# a_n945_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X20 a_15_n75# a_n1167_n101# a_n81_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X21 a_n81_n75# a_n1167_n101# a_n177_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X22 a_111_n75# a_n1167_n101# a_15_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X23 a_n273_n75# a_n1167_n101# a_n369_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X24 a_n177_n75# a_n1167_n101# a_n273_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
C0 a_399_n75# a_687_n75# 0.05fF
C1 a_n369_n75# a_n753_n75# 0.03fF
C2 a_1167_n75# a_879_n75# 0.05fF
C3 a_15_n75# a_303_n75# 0.05fF
C4 a_n369_n75# a_n657_n75# 0.05fF
C5 a_207_n75# a_495_n75# 0.05fF
C6 a_15_n75# a_399_n75# 0.03fF
C7 a_n177_n75# a_111_n75# 0.05fF
C8 a_n465_n75# a_n561_n75# 0.22fF
C9 a_591_n75# a_783_n75# 0.08fF
C10 a_879_n75# a_687_n75# 0.08fF
C11 a_n465_n75# a_n753_n75# 0.05fF
C12 a_n1229_n75# a_n945_n75# 0.05fF
C13 a_n273_n75# a_n561_n75# 0.05fF
C14 a_975_n75# a_879_n75# 0.22fF
C15 a_n465_n75# a_n657_n75# 0.08fF
C16 a_15_n75# a_n177_n75# 0.08fF
C17 a_n1137_n75# a_n1041_n75# 0.22fF
C18 a_591_n75# a_495_n75# 0.22fF
C19 a_n561_n75# a_n849_n75# 0.05fF
C20 a_111_n75# a_n81_n75# 0.08fF
C21 a_207_n75# a_111_n75# 0.22fF
C22 a_n273_n75# a_n657_n75# 0.03fF
C23 a_n753_n75# a_n849_n75# 0.22fF
C24 a_399_n75# a_303_n75# 0.22fF
C25 a_n657_n75# a_n849_n75# 0.08fF
C26 a_n945_n75# a_n849_n75# 0.22fF
C27 a_15_n75# a_n369_n75# 0.03fF
C28 a_15_n75# a_n81_n75# 0.22fF
C29 a_15_n75# a_207_n75# 0.08fF
C30 a_1071_n75# a_879_n75# 0.08fF
C31 a_n273_n75# a_111_n75# 0.03fF
C32 a_495_n75# a_783_n75# 0.05fF
C33 a_n561_n75# a_n753_n75# 0.08fF
C34 a_591_n75# a_687_n75# 0.22fF
C35 a_n657_n75# a_n561_n75# 0.22fF
C36 a_n945_n75# a_n561_n75# 0.03fF
C37 a_591_n75# a_975_n75# 0.03fF
C38 a_15_n75# a_n273_n75# 0.05fF
C39 a_n1229_n75# a_n1041_n75# 0.08fF
C40 a_n945_n75# a_n753_n75# 0.08fF
C41 a_n657_n75# a_n753_n75# 0.22fF
C42 a_1167_n75# a_783_n75# 0.03fF
C43 a_n945_n75# a_n657_n75# 0.05fF
C44 a_303_n75# a_n81_n75# 0.03fF
C45 a_207_n75# a_303_n75# 0.22fF
C46 a_399_n75# a_207_n75# 0.08fF
C47 a_687_n75# a_783_n75# 0.22fF
C48 a_n849_n75# a_n1041_n75# 0.08fF
C49 a_975_n75# a_783_n75# 0.08fF
C50 a_495_n75# a_111_n75# 0.03fF
C51 a_n177_n75# a_n369_n75# 0.08fF
C52 a_591_n75# a_303_n75# 0.05fF
C53 a_n177_n75# a_n81_n75# 0.22fF
C54 a_495_n75# a_687_n75# 0.08fF
C55 a_n1137_n75# a_n1229_n75# 0.22fF
C56 a_207_n75# a_n177_n75# 0.03fF
C57 a_399_n75# a_591_n75# 0.08fF
C58 a_n465_n75# a_n177_n75# 0.05fF
C59 a_n369_n75# a_n81_n75# 0.05fF
C60 a_n753_n75# a_n1041_n75# 0.05fF
C61 a_n1137_n75# a_n849_n75# 0.05fF
C62 a_207_n75# a_n81_n75# 0.05fF
C63 a_591_n75# a_879_n75# 0.05fF
C64 a_1167_n75# a_975_n75# 0.08fF
C65 a_1071_n75# a_783_n75# 0.05fF
C66 a_n273_n75# a_n177_n75# 0.22fF
C67 a_n945_n75# a_n1041_n75# 0.22fF
C68 a_n657_n75# a_n1041_n75# 0.03fF
C69 a_n465_n75# a_n369_n75# 0.22fF
C70 a_399_n75# a_783_n75# 0.03fF
C71 a_15_n75# a_111_n75# 0.22fF
C72 a_n465_n75# a_n81_n75# 0.03fF
C73 a_975_n75# a_687_n75# 0.05fF
C74 a_n273_n75# a_n369_n75# 0.22fF
C75 a_303_n75# a_495_n75# 0.08fF
C76 a_207_n75# a_591_n75# 0.03fF
C77 a_n273_n75# a_n81_n75# 0.08fF
C78 a_399_n75# a_495_n75# 0.22fF
C79 a_879_n75# a_783_n75# 0.22fF
C80 a_n1137_n75# a_n753_n75# 0.03fF
C81 a_1167_n75# a_1071_n75# 0.22fF
C82 a_n177_n75# a_n561_n75# 0.03fF
C83 a_n1137_n75# a_n945_n75# 0.08fF
C84 a_n465_n75# a_n273_n75# 0.08fF
C85 a_495_n75# a_879_n75# 0.03fF
C86 a_n1229_n75# a_n849_n75# 0.03fF
C87 a_303_n75# a_111_n75# 0.08fF
C88 a_n465_n75# a_n849_n75# 0.03fF
C89 a_1071_n75# a_687_n75# 0.03fF
C90 a_399_n75# a_111_n75# 0.05fF
C91 a_n369_n75# a_n561_n75# 0.08fF
C92 a_1071_n75# a_975_n75# 0.22fF
C93 a_303_n75# a_687_n75# 0.03fF
C94 a_1167_n75# w_n1367_n285# 0.10fF
C95 a_1071_n75# w_n1367_n285# 0.07fF
C96 a_975_n75# w_n1367_n285# 0.06fF
C97 a_879_n75# w_n1367_n285# 0.05fF
C98 a_783_n75# w_n1367_n285# 0.04fF
C99 a_687_n75# w_n1367_n285# 0.04fF
C100 a_591_n75# w_n1367_n285# 0.04fF
C101 a_495_n75# w_n1367_n285# 0.04fF
C102 a_399_n75# w_n1367_n285# 0.04fF
C103 a_303_n75# w_n1367_n285# 0.04fF
C104 a_207_n75# w_n1367_n285# 0.04fF
C105 a_111_n75# w_n1367_n285# 0.04fF
C106 a_15_n75# w_n1367_n285# 0.04fF
C107 a_n81_n75# w_n1367_n285# 0.04fF
C108 a_n177_n75# w_n1367_n285# 0.04fF
C109 a_n273_n75# w_n1367_n285# 0.04fF
C110 a_n369_n75# w_n1367_n285# 0.04fF
C111 a_n465_n75# w_n1367_n285# 0.04fF
C112 a_n561_n75# w_n1367_n285# 0.04fF
C113 a_n657_n75# w_n1367_n285# 0.04fF
C114 a_n753_n75# w_n1367_n285# 0.04fF
C115 a_n849_n75# w_n1367_n285# 0.04fF
C116 a_n945_n75# w_n1367_n285# 0.04fF
C117 a_n1041_n75# w_n1367_n285# 0.04fF
C118 a_n1137_n75# w_n1367_n285# 0.04fF
C119 a_n1229_n75# w_n1367_n285# 0.04fF
C120 a_n1167_n101# w_n1367_n285# 2.55fF
.ends

.subckt sky130_fd_pr__nfet_01v8_MUHGM9 a_33_n101# a_n129_n75# a_735_n75# a_255_n75#
+ a_n417_n75# a_n989_n75# a_63_n75# a_543_n75# a_n705_n75# a_n225_n75# a_n33_n75#
+ a_831_n75# a_351_n75# a_n927_n101# a_n513_n75# a_n897_n75# w_n1127_n285# a_639_n75#
+ a_159_n75# a_n801_n75# a_n321_n75# a_927_n75# a_447_n75# a_n609_n75#
X0 a_63_n75# a_33_n101# a_n33_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_927_n75# a_33_n101# a_831_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_n33_n75# a_n927_n101# a_n129_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_159_n75# a_33_n101# a_63_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_255_n75# a_33_n101# a_159_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_351_n75# a_33_n101# a_255_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_447_n75# a_33_n101# a_351_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_543_n75# a_33_n101# a_447_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_735_n75# a_33_n101# a_639_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_831_n75# a_33_n101# a_735_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_639_n75# a_33_n101# a_543_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n321_n75# a_n927_n101# a_n417_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_n801_n75# a_n927_n101# a_n897_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n705_n75# a_n927_n101# a_n801_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n513_n75# a_n927_n101# a_n609_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n417_n75# a_n927_n101# a_n513_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n225_n75# a_n927_n101# a_n321_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n129_n75# a_n927_n101# a_n225_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_n897_n75# a_n927_n101# a_n989_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n609_n75# a_n927_n101# a_n705_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
C0 a_159_n75# a_447_n75# 0.05fF
C1 a_n705_n75# a_n989_n75# 0.05fF
C2 a_n705_n75# a_n513_n75# 0.08fF
C3 a_n321_n75# a_n33_n75# 0.05fF
C4 a_831_n75# a_543_n75# 0.05fF
C5 a_n609_n75# a_n417_n75# 0.08fF
C6 a_n321_n75# a_63_n75# 0.03fF
C7 a_n513_n75# a_n225_n75# 0.05fF
C8 a_735_n75# a_639_n75# 0.22fF
C9 a_n33_n75# a_255_n75# 0.05fF
C10 a_63_n75# a_255_n75# 0.08fF
C11 a_n705_n75# a_n417_n75# 0.05fF
C12 a_n897_n75# a_n989_n75# 0.22fF
C13 a_n513_n75# a_n897_n75# 0.03fF
C14 a_735_n75# a_351_n75# 0.03fF
C15 a_735_n75# a_543_n75# 0.08fF
C16 a_n321_n75# a_n513_n75# 0.08fF
C17 a_639_n75# a_447_n75# 0.08fF
C18 a_n225_n75# a_n417_n75# 0.08fF
C19 a_n129_n75# a_n225_n75# 0.22fF
C20 a_351_n75# a_159_n75# 0.08fF
C21 a_159_n75# a_543_n75# 0.03fF
C22 a_63_n75# a_n33_n75# 0.22fF
C23 a_351_n75# a_447_n75# 0.22fF
C24 a_543_n75# a_447_n75# 0.22fF
C25 a_n321_n75# a_n417_n75# 0.22fF
C26 a_n321_n75# a_n129_n75# 0.08fF
C27 a_n801_n75# a_n989_n75# 0.08fF
C28 a_n513_n75# a_n801_n75# 0.05fF
C29 a_159_n75# a_n225_n75# 0.03fF
C30 a_n129_n75# a_255_n75# 0.03fF
C31 a_351_n75# a_639_n75# 0.05fF
C32 a_543_n75# a_639_n75# 0.22fF
C33 a_n801_n75# a_n417_n75# 0.03fF
C34 a_351_n75# a_543_n75# 0.08fF
C35 a_n33_n75# a_n417_n75# 0.03fF
C36 a_n129_n75# a_n33_n75# 0.22fF
C37 a_159_n75# a_255_n75# 0.22fF
C38 a_63_n75# a_n129_n75# 0.08fF
C39 a_n705_n75# a_n609_n75# 0.22fF
C40 a_927_n75# a_831_n75# 0.22fF
C41 a_n927_n101# a_33_n101# 0.08fF
C42 a_447_n75# a_255_n75# 0.08fF
C43 a_n609_n75# a_n225_n75# 0.03fF
C44 a_n513_n75# a_n417_n75# 0.22fF
C45 a_n129_n75# a_n513_n75# 0.03fF
C46 a_159_n75# a_n33_n75# 0.08fF
C47 a_735_n75# a_927_n75# 0.08fF
C48 a_n897_n75# a_n609_n75# 0.05fF
C49 a_63_n75# a_159_n75# 0.22fF
C50 a_n321_n75# a_n609_n75# 0.05fF
C51 a_639_n75# a_255_n75# 0.03fF
C52 a_63_n75# a_447_n75# 0.03fF
C53 a_n129_n75# a_n417_n75# 0.05fF
C54 a_n705_n75# a_n897_n75# 0.08fF
C55 a_351_n75# a_255_n75# 0.22fF
C56 a_543_n75# a_255_n75# 0.05fF
C57 a_n321_n75# a_n705_n75# 0.03fF
C58 a_735_n75# a_831_n75# 0.22fF
C59 a_n321_n75# a_n225_n75# 0.22fF
C60 a_n801_n75# a_n609_n75# 0.08fF
C61 a_927_n75# a_639_n75# 0.05fF
C62 a_351_n75# a_n33_n75# 0.03fF
C63 a_n129_n75# a_159_n75# 0.05fF
C64 a_831_n75# a_447_n75# 0.03fF
C65 a_63_n75# a_351_n75# 0.05fF
C66 a_n705_n75# a_n801_n75# 0.22fF
C67 a_927_n75# a_543_n75# 0.03fF
C68 a_n609_n75# a_n989_n75# 0.03fF
C69 a_n513_n75# a_n609_n75# 0.22fF
C70 a_n33_n75# a_n225_n75# 0.08fF
C71 a_735_n75# a_447_n75# 0.05fF
C72 a_63_n75# a_n225_n75# 0.05fF
C73 a_831_n75# a_639_n75# 0.08fF
C74 a_n801_n75# a_n897_n75# 0.22fF
C75 a_927_n75# w_n1127_n285# 0.04fF
C76 a_831_n75# w_n1127_n285# 0.04fF
C77 a_735_n75# w_n1127_n285# 0.04fF
C78 a_639_n75# w_n1127_n285# 0.04fF
C79 a_543_n75# w_n1127_n285# 0.04fF
C80 a_447_n75# w_n1127_n285# 0.04fF
C81 a_351_n75# w_n1127_n285# 0.04fF
C82 a_255_n75# w_n1127_n285# 0.04fF
C83 a_159_n75# w_n1127_n285# 0.04fF
C84 a_63_n75# w_n1127_n285# 0.04fF
C85 a_n33_n75# w_n1127_n285# 0.04fF
C86 a_n129_n75# w_n1127_n285# 0.04fF
C87 a_n225_n75# w_n1127_n285# 0.04fF
C88 a_n321_n75# w_n1127_n285# 0.04fF
C89 a_n417_n75# w_n1127_n285# 0.04fF
C90 a_n513_n75# w_n1127_n285# 0.04fF
C91 a_n609_n75# w_n1127_n285# 0.04fF
C92 a_n705_n75# w_n1127_n285# 0.04fF
C93 a_n801_n75# w_n1127_n285# 0.04fF
C94 a_n897_n75# w_n1127_n285# 0.04fF
C95 a_n989_n75# w_n1127_n285# 0.04fF
C96 a_33_n101# w_n1127_n285# 0.99fF
C97 a_n927_n101# w_n1127_n285# 0.99fF
.ends

.subckt sky130_fd_pr__pfet_01v8_NKZXKB VSUBS a_33_n247# a_n801_n150# a_n417_n150#
+ a_351_n150# a_255_n150# a_n705_n150# a_n609_n150# a_159_n150# a_543_n150# a_447_n150#
+ a_831_n150# a_n897_n150# a_n33_n150# a_735_n150# a_n927_n247# a_639_n150# a_n321_n150#
+ a_927_n150# a_n225_n150# a_63_n150# a_n989_n150# a_n513_n150# a_n129_n150# w_n1127_n369#
X0 a_n513_n150# a_n927_n247# a_n609_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_63_n150# a_33_n247# a_n33_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_735_n150# a_33_n247# a_639_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n801_n150# a_n927_n247# a_n897_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n927_n247# a_n225_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n927_n247# a_n513_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_639_n150# a_33_n247# a_543_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n705_n150# a_n927_n247# a_n801_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n33_n150# a_n927_n247# a_n129_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_351_n150# a_33_n247# a_255_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_n609_n150# a_n927_n247# a_n705_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n897_n150# a_n927_n247# a_n989_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_927_n150# a_33_n247# a_831_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_255_n150# a_33_n247# a_159_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n321_n150# a_n927_n247# a_n417_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_543_n150# a_33_n247# a_447_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_831_n150# a_33_n247# a_735_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_159_n150# a_33_n247# a_63_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_n225_n150# a_n927_n247# a_n321_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_447_n150# a_33_n247# a_351_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n989_n150# a_n609_n150# 0.07fF
C1 a_447_n150# a_159_n150# 0.10fF
C2 a_447_n150# a_639_n150# 0.16fF
C3 a_543_n150# a_735_n150# 0.16fF
C4 a_63_n150# a_n321_n150# 0.07fF
C5 a_n513_n150# a_n897_n150# 0.07fF
C6 a_n417_n150# a_n129_n150# 0.10fF
C7 a_927_n150# a_831_n150# 0.43fF
C8 a_n321_n150# a_n129_n150# 0.16fF
C9 a_447_n150# a_735_n150# 0.10fF
C10 a_255_n150# a_159_n150# 0.43fF
C11 a_639_n150# a_255_n150# 0.07fF
C12 a_n801_n150# a_n897_n150# 0.43fF
C13 a_63_n150# a_159_n150# 0.43fF
C14 a_927_n150# a_543_n150# 0.07fF
C15 a_n513_n150# a_n609_n150# 0.43fF
C16 a_n33_n150# a_n225_n150# 0.16fF
C17 a_159_n150# a_n129_n150# 0.10fF
C18 a_n321_n150# a_n417_n150# 0.43fF
C19 a_n801_n150# a_n609_n150# 0.16fF
C20 a_n897_n150# a_n705_n150# 0.16fF
C21 a_351_n150# a_159_n150# 0.16fF
C22 a_639_n150# a_351_n150# 0.10fF
C23 a_n225_n150# a_n609_n150# 0.07fF
C24 a_543_n150# a_831_n150# 0.10fF
C25 a_n513_n150# a_n129_n150# 0.07fF
C26 a_n609_n150# a_n705_n150# 0.43fF
C27 a_63_n150# a_n225_n150# 0.10fF
C28 a_351_n150# a_735_n150# 0.07fF
C29 a_447_n150# a_831_n150# 0.07fF
C30 a_n513_n150# a_n417_n150# 0.43fF
C31 a_n225_n150# a_n129_n150# 0.43fF
C32 a_n321_n150# a_n513_n150# 0.16fF
C33 a_447_n150# a_543_n150# 0.43fF
C34 a_n801_n150# a_n417_n150# 0.07fF
C35 a_639_n150# a_735_n150# 0.43fF
C36 a_n989_n150# a_n801_n150# 0.16fF
C37 a_n897_n150# a_n609_n150# 0.10fF
C38 a_n225_n150# a_n417_n150# 0.16fF
C39 a_255_n150# a_543_n150# 0.10fF
C40 a_n321_n150# a_n225_n150# 0.43fF
C41 a_n33_n150# a_255_n150# 0.10fF
C42 a_n417_n150# a_n705_n150# 0.10fF
C43 a_63_n150# a_n33_n150# 0.43fF
C44 a_n321_n150# a_n705_n150# 0.07fF
C45 a_n989_n150# a_n705_n150# 0.10fF
C46 a_447_n150# a_255_n150# 0.16fF
C47 a_927_n150# a_639_n150# 0.10fF
C48 a_n225_n150# a_159_n150# 0.07fF
C49 a_n33_n150# a_n129_n150# 0.43fF
C50 a_63_n150# a_447_n150# 0.07fF
C51 a_n927_n247# a_33_n247# 0.09fF
C52 a_n513_n150# a_n801_n150# 0.10fF
C53 a_351_n150# a_543_n150# 0.16fF
C54 a_n33_n150# a_351_n150# 0.07fF
C55 a_927_n150# a_735_n150# 0.16fF
C56 a_n33_n150# a_n417_n150# 0.07fF
C57 a_n513_n150# a_n225_n150# 0.10fF
C58 a_63_n150# a_255_n150# 0.16fF
C59 a_n321_n150# a_n33_n150# 0.10fF
C60 a_447_n150# a_351_n150# 0.43fF
C61 a_639_n150# a_831_n150# 0.16fF
C62 a_n513_n150# a_n705_n150# 0.16fF
C63 a_255_n150# a_n129_n150# 0.07fF
C64 a_n989_n150# a_n897_n150# 0.43fF
C65 a_63_n150# a_n129_n150# 0.16fF
C66 a_543_n150# a_159_n150# 0.07fF
C67 a_639_n150# a_543_n150# 0.43fF
C68 a_n801_n150# a_n705_n150# 0.43fF
C69 a_n417_n150# a_n609_n150# 0.16fF
C70 a_n33_n150# a_159_n150# 0.16fF
C71 a_n321_n150# a_n609_n150# 0.10fF
C72 a_735_n150# a_831_n150# 0.43fF
C73 a_351_n150# a_255_n150# 0.43fF
C74 a_63_n150# a_351_n150# 0.10fF
C75 a_927_n150# VSUBS 0.03fF
C76 a_831_n150# VSUBS 0.03fF
C77 a_735_n150# VSUBS 0.03fF
C78 a_639_n150# VSUBS 0.03fF
C79 a_543_n150# VSUBS 0.03fF
C80 a_447_n150# VSUBS 0.03fF
C81 a_351_n150# VSUBS 0.03fF
C82 a_255_n150# VSUBS 0.03fF
C83 a_159_n150# VSUBS 0.03fF
C84 a_63_n150# VSUBS 0.03fF
C85 a_n33_n150# VSUBS 0.03fF
C86 a_n129_n150# VSUBS 0.03fF
C87 a_n225_n150# VSUBS 0.03fF
C88 a_n321_n150# VSUBS 0.03fF
C89 a_n417_n150# VSUBS 0.03fF
C90 a_n513_n150# VSUBS 0.03fF
C91 a_n609_n150# VSUBS 0.03fF
C92 a_n705_n150# VSUBS 0.03fF
C93 a_n801_n150# VSUBS 0.03fF
C94 a_n897_n150# VSUBS 0.03fF
C95 a_n989_n150# VSUBS 0.03fF
C96 a_33_n247# VSUBS 1.04fF
C97 a_n927_n247# VSUBS 1.04fF
C98 w_n1127_n369# VSUBS 6.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_8GRULZ a_n1761_n132# a_1045_n44# a_n1461_n44# a_n1103_n44#
+ a_n29_n44# a_n387_n44# a_1761_n44# a_n1819_n44# a_1403_n44# a_687_n44# w_n1957_n254#
+ a_329_n44# a_n745_n44#
X0 a_329_n44# a_n1761_n132# a_n29_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X1 a_1761_n44# a_n1761_n132# a_1403_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X2 a_n745_n44# a_n1761_n132# a_n1103_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X3 a_1045_n44# a_n1761_n132# a_687_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X4 a_n29_n44# a_n1761_n132# a_n387_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X5 a_n1103_n44# a_n1761_n132# a_n1461_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X6 a_n387_n44# a_n1761_n132# a_n745_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X7 a_687_n44# a_n1761_n132# a_329_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X8 a_1403_n44# a_n1761_n132# a_1045_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X9 a_n1461_n44# a_n1761_n132# a_n1819_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
C0 a_n745_n44# a_n1103_n44# 0.04fF
C1 a_329_n44# a_n29_n44# 0.04fF
C2 a_n745_n44# a_n387_n44# 0.04fF
C3 a_687_n44# a_1045_n44# 0.04fF
C4 a_n1819_n44# a_n1461_n44# 0.04fF
C5 a_329_n44# a_687_n44# 0.04fF
C6 a_1761_n44# a_1403_n44# 0.04fF
C7 a_1403_n44# a_1045_n44# 0.04fF
C8 a_n29_n44# a_n387_n44# 0.04fF
C9 a_n1461_n44# a_n1103_n44# 0.04fF
C10 a_1761_n44# w_n1957_n254# 0.04fF
C11 a_1403_n44# w_n1957_n254# 0.04fF
C12 a_1045_n44# w_n1957_n254# 0.04fF
C13 a_687_n44# w_n1957_n254# 0.04fF
C14 a_329_n44# w_n1957_n254# 0.04fF
C15 a_n29_n44# w_n1957_n254# 0.04fF
C16 a_n387_n44# w_n1957_n254# 0.04fF
C17 a_n745_n44# w_n1957_n254# 0.04fF
C18 a_n1103_n44# w_n1957_n254# 0.04fF
C19 a_n1461_n44# w_n1957_n254# 0.04fF
C20 a_n1819_n44# w_n1957_n254# 0.04fF
C21 a_n1761_n132# w_n1957_n254# 3.23fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ND88ZC VSUBS a_303_n150# a_n753_n150# a_n369_n150#
+ w_n1367_n369# a_207_n150# a_n657_n150# a_591_n150# a_n1229_n150# a_n945_n150# a_495_n150#
+ a_n1041_n150# a_n849_n150# a_n81_n150# a_399_n150# a_783_n150# a_1071_n150# a_687_n150#
+ a_975_n150# a_n1137_n150# a_n273_n150# a_111_n150# a_879_n150# a_n177_n150# a_n561_n150#
+ a_15_n150# a_1167_n150# a_n1167_n247# a_n465_n150#
X0 a_n1137_n150# a_n1167_n247# a_n1229_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_495_n150# a_n1167_n247# a_399_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n561_n150# a_n1167_n247# a_n657_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_111_n150# a_n1167_n247# a_15_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_783_n150# a_n1167_n247# a_687_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_1071_n150# a_n1167_n247# a_975_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_399_n150# a_n1167_n247# a_303_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n465_n150# a_n1167_n247# a_n561_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_687_n150# a_n1167_n247# a_591_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n753_n150# a_n1167_n247# a_n849_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_975_n150# a_n1167_n247# a_879_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n81_n150# a_n1167_n247# a_n177_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_15_n150# a_n1167_n247# a_n81_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_n1041_n150# a_n1167_n247# a_n1137_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n369_n150# a_n1167_n247# a_n465_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_n657_n150# a_n1167_n247# a_n753_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_879_n150# a_n1167_n247# a_783_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_n945_n150# a_n1167_n247# a_n1041_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_1167_n150# a_n1167_n247# a_1071_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_303_n150# a_n1167_n247# a_207_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X20 a_n273_n150# a_n1167_n247# a_n369_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X21 a_591_n150# a_n1167_n247# a_495_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X22 a_n849_n150# a_n1167_n247# a_n945_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_207_n150# a_n1167_n247# a_111_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X24 a_n177_n150# a_n1167_n247# a_n273_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n657_n150# a_n273_n150# 0.07fF
C1 a_n849_n150# a_n945_n150# 0.43fF
C2 a_687_n150# a_1071_n150# 0.07fF
C3 a_783_n150# a_687_n150# 0.43fF
C4 a_n1137_n150# a_n849_n150# 0.10fF
C5 a_n81_n150# a_111_n150# 0.16fF
C6 a_n753_n150# a_n561_n150# 0.16fF
C7 a_n657_n150# a_n945_n150# 0.10fF
C8 a_n177_n150# a_n561_n150# 0.07fF
C9 a_207_n150# a_111_n150# 0.43fF
C10 a_687_n150# a_303_n150# 0.07fF
C11 a_207_n150# a_591_n150# 0.07fF
C12 a_n945_n150# a_n1041_n150# 0.43fF
C13 a_n465_n150# a_n561_n150# 0.43fF
C14 a_n1137_n150# a_n1041_n150# 0.43fF
C15 a_1167_n150# a_975_n150# 0.16fF
C16 w_n1367_n369# a_975_n150# 0.05fF
C17 a_1167_n150# a_879_n150# 0.10fF
C18 w_n1367_n369# a_879_n150# 0.04fF
C19 a_n273_n150# a_15_n150# 0.10fF
C20 a_207_n150# a_495_n150# 0.10fF
C21 a_n177_n150# a_n273_n150# 0.43fF
C22 a_303_n150# a_15_n150# 0.10fF
C23 a_n753_n150# a_n945_n150# 0.16fF
C24 a_n465_n150# a_n273_n150# 0.16fF
C25 a_n1137_n150# a_n753_n150# 0.07fF
C26 a_n81_n150# a_n273_n150# 0.16fF
C27 a_n561_n150# a_n369_n150# 0.16fF
C28 a_1167_n150# a_1071_n150# 0.43fF
C29 a_783_n150# a_1167_n150# 0.07fF
C30 w_n1367_n369# a_1071_n150# 0.07fF
C31 a_n657_n150# a_n849_n150# 0.16fF
C32 a_n81_n150# a_303_n150# 0.07fF
C33 a_687_n150# a_399_n150# 0.10fF
C34 a_n849_n150# a_n1041_n150# 0.16fF
C35 a_591_n150# a_975_n150# 0.07fF
C36 a_207_n150# a_303_n150# 0.43fF
C37 a_495_n150# a_111_n150# 0.07fF
C38 a_879_n150# a_591_n150# 0.10fF
C39 a_n273_n150# a_n369_n150# 0.43fF
C40 a_495_n150# a_591_n150# 0.43fF
C41 a_879_n150# a_975_n150# 0.43fF
C42 a_n657_n150# a_n1041_n150# 0.07fF
C43 a_399_n150# a_15_n150# 0.07fF
C44 a_495_n150# a_879_n150# 0.07fF
C45 a_n849_n150# a_n753_n150# 0.43fF
C46 a_783_n150# a_591_n150# 0.16fF
C47 a_n273_n150# a_111_n150# 0.07fF
C48 a_1071_n150# a_975_n150# 0.43fF
C49 a_783_n150# a_975_n150# 0.16fF
C50 a_879_n150# a_1071_n150# 0.16fF
C51 a_783_n150# a_879_n150# 0.43fF
C52 a_n657_n150# a_n753_n150# 0.43fF
C53 a_303_n150# a_111_n150# 0.16fF
C54 a_783_n150# a_495_n150# 0.10fF
C55 a_n465_n150# a_n849_n150# 0.07fF
C56 a_591_n150# a_303_n150# 0.10fF
C57 a_207_n150# a_399_n150# 0.16fF
C58 a_n753_n150# a_n1041_n150# 0.10fF
C59 a_783_n150# a_1071_n150# 0.10fF
C60 a_n657_n150# a_n465_n150# 0.16fF
C61 a_n561_n150# a_n273_n150# 0.10fF
C62 a_495_n150# a_303_n150# 0.16fF
C63 a_n1229_n150# a_n945_n150# 0.10fF
C64 a_n1137_n150# a_n1229_n150# 0.43fF
C65 a_n945_n150# a_n561_n150# 0.07fF
C66 a_n657_n150# a_n369_n150# 0.10fF
C67 a_n177_n150# a_15_n150# 0.16fF
C68 a_399_n150# a_111_n150# 0.10fF
C69 a_399_n150# a_591_n150# 0.16fF
C70 a_n465_n150# a_n753_n150# 0.10fF
C71 a_n177_n150# a_n465_n150# 0.10fF
C72 a_n81_n150# a_15_n150# 0.43fF
C73 a_n81_n150# a_n177_n150# 0.43fF
C74 a_399_n150# a_495_n150# 0.43fF
C75 a_207_n150# a_15_n150# 0.16fF
C76 a_n177_n150# a_207_n150# 0.07fF
C77 a_n1229_n150# a_n849_n150# 0.07fF
C78 a_n1137_n150# a_n945_n150# 0.16fF
C79 a_n81_n150# a_n465_n150# 0.07fF
C80 a_n849_n150# a_n561_n150# 0.10fF
C81 a_n753_n150# a_n369_n150# 0.07fF
C82 a_783_n150# a_399_n150# 0.07fF
C83 a_15_n150# a_n369_n150# 0.07fF
C84 a_n177_n150# a_n369_n150# 0.16fF
C85 a_687_n150# a_591_n150# 0.43fF
C86 a_n81_n150# a_207_n150# 0.10fF
C87 a_n657_n150# a_n561_n150# 0.43fF
C88 a_687_n150# a_975_n150# 0.10fF
C89 a_687_n150# a_879_n150# 0.16fF
C90 a_n465_n150# a_n369_n150# 0.43fF
C91 a_n1229_n150# a_n1041_n150# 0.16fF
C92 a_399_n150# a_303_n150# 0.43fF
C93 a_n81_n150# a_n369_n150# 0.10fF
C94 a_687_n150# a_495_n150# 0.16fF
C95 a_1167_n150# w_n1367_n369# 0.14fF
C96 a_15_n150# a_111_n150# 0.43fF
C97 a_n177_n150# a_111_n150# 0.10fF
C98 a_1167_n150# VSUBS 0.03fF
C99 a_1071_n150# VSUBS 0.03fF
C100 a_975_n150# VSUBS 0.03fF
C101 a_879_n150# VSUBS 0.03fF
C102 a_783_n150# VSUBS 0.03fF
C103 a_687_n150# VSUBS 0.03fF
C104 a_591_n150# VSUBS 0.03fF
C105 a_495_n150# VSUBS 0.03fF
C106 a_399_n150# VSUBS 0.03fF
C107 a_303_n150# VSUBS 0.03fF
C108 a_207_n150# VSUBS 0.03fF
C109 a_111_n150# VSUBS 0.03fF
C110 a_15_n150# VSUBS 0.03fF
C111 a_n81_n150# VSUBS 0.03fF
C112 a_n177_n150# VSUBS 0.03fF
C113 a_n273_n150# VSUBS 0.03fF
C114 a_n369_n150# VSUBS 0.03fF
C115 a_n465_n150# VSUBS 0.03fF
C116 a_n561_n150# VSUBS 0.03fF
C117 a_n657_n150# VSUBS 0.03fF
C118 a_n753_n150# VSUBS 0.03fF
C119 a_n849_n150# VSUBS 0.03fF
C120 a_n945_n150# VSUBS 0.03fF
C121 a_n1041_n150# VSUBS 0.03fF
C122 a_n1137_n150# VSUBS 0.03fF
C123 a_n1229_n150# VSUBS 0.03fF
C124 a_n1167_n247# VSUBS 2.63fF
C125 w_n1367_n369# VSUBS 7.85fF
.ends

.subckt charge_pump nswitch vss vdd nUp Down w_2544_775# out pswitch iref nDown biasp
+ Up w_6648_570#
Xsky130_fd_pr__pfet_01v8_4ML9WA_0 vss pswitch vdd pswitch pswitch pswitch nUp pswitch
+ pswitch pswitch pswitch pswitch pswitch pswitch sky130_fd_pr__pfet_01v8_4ML9WA
Xsky130_fd_pr__nfet_01v8_YCGG98_0 vss out out vss vss vss out out vss vss out vss
+ out out out vss out vss out out out vss vss vss out vss vss nswitch sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_1 iref vss vss iref iref iref vss vss iref iref vss
+ iref vss vss vss iref vss iref vss vss vss vss iref iref vss iref iref iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_2 biasp vss vss biasp biasp biasp vss vss biasp biasp
+ vss biasp vss vss vss biasp vss biasp vss vss vss vss biasp biasp vss biasp biasp
+ iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_MUHGM9_0 nDown iref nswitch vss nswitch nswitch vss nswitch
+ iref nswitch nswitch vss nswitch Down iref iref vss vss nswitch nswitch iref nswitch
+ vss nswitch sky130_fd_pr__nfet_01v8_MUHGM9
Xsky130_fd_pr__pfet_01v8_NKZXKB_0 vss Up pswitch pswitch pswitch vdd biasp pswitch
+ pswitch pswitch vdd vdd biasp pswitch pswitch nUp vdd biasp pswitch pswitch vdd
+ pswitch biasp biasp vdd sky130_fd_pr__pfet_01v8_NKZXKB
Xsky130_fd_pr__nfet_01v8_8GRULZ_0 Down nswitch nswitch nswitch nswitch nswitch nswitch
+ nswitch nswitch nswitch vss nswitch nswitch sky130_fd_pr__nfet_01v8_8GRULZ
Xsky130_fd_pr__pfet_01v8_ND88ZC_0 vss vdd out out vdd out vdd out vdd out vdd vdd
+ vdd vdd out out vdd vdd out out vdd vdd vdd out out out out pswitch vdd sky130_fd_pr__pfet_01v8_ND88ZC
Xsky130_fd_pr__pfet_01v8_ND88ZC_1 vss biasp vdd vdd vdd vdd biasp vdd biasp vdd biasp
+ biasp biasp biasp vdd vdd biasp biasp vdd vdd biasp biasp biasp vdd vdd vdd vdd
+ biasp biasp sky130_fd_pr__pfet_01v8_ND88ZC
C0 pswitch biasp 3.11fF
C1 vdd pswitch 3.98fF
C2 nDown Down 0.13fF
C3 iref biasp 0.80fF
C4 pswitch nswitch 0.06fF
C5 iref nswitch 1.91fF
C6 nUp pswitch 5.66fF
C7 out vdd 6.66fF
C8 nDown nswitch 0.31fF
C9 out nswitch 1.28fF
C10 Down nswitch 2.27fF
C11 vdd biasp 2.64fF
C12 out pswitch 4.91fF
C13 pswitch Up 0.70fF
C14 biasp nswitch 0.03fF
C15 nUp out 0.31fF
C16 nUp Down 0.25fF
C17 nUp Up 0.15fF
C18 vdd nswitch 0.07fF
C19 vdd vss 35.71fF
C20 Down vss 4.77fF
C21 Up vss 1.17fF
C22 nswitch vss 6.39fF
C23 nDown vss 1.11fF
C24 biasp vss 8.73fF
C25 iref vss 10.12fF
C26 out vss -3.49fF
C27 pswitch vss 3.45fF
C28 nUp vss 5.85fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MACBVW VSUBS m3_n2650_n13200# m3_n7969_n2600# m3_7988_8000#
+ m3_2669_n7900# m3_n13288_n2600# m3_n2650_2700# m3_2669_2700# m3_n13288_n13200# m3_n7969_n13200#
+ m3_n13288_8000# m3_7988_2700# m3_n2650_n7900# m3_7988_n7900# m3_2669_n13200# m3_n7969_8000#
+ m3_n13288_2700# m3_n7969_n7900# m3_n13288_n7900# m3_2669_n2600# m3_n7969_2700# m3_7988_n13200#
+ c1_n13188_n13100# m3_7988_n2600# m3_n2650_n2600# m3_n2650_8000# m3_2669_8000#
X0 c1_n13188_n13100# m3_2669_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X1 c1_n13188_n13100# m3_n2650_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X2 c1_n13188_n13100# m3_2669_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X3 c1_n13188_n13100# m3_n13288_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X4 c1_n13188_n13100# m3_n7969_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X5 c1_n13188_n13100# m3_n13288_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X6 c1_n13188_n13100# m3_2669_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X7 c1_n13188_n13100# m3_7988_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X8 c1_n13188_n13100# m3_2669_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X9 c1_n13188_n13100# m3_7988_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X10 c1_n13188_n13100# m3_n7969_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X11 c1_n13188_n13100# m3_7988_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X12 c1_n13188_n13100# m3_n7969_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X13 c1_n13188_n13100# m3_7988_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X14 c1_n13188_n13100# m3_n13288_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X15 c1_n13188_n13100# m3_n7969_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X16 c1_n13188_n13100# m3_n2650_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X17 c1_n13188_n13100# m3_n2650_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X18 c1_n13188_n13100# m3_n2650_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X19 c1_n13188_n13100# m3_7988_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X20 c1_n13188_n13100# m3_n13288_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X21 c1_n13188_n13100# m3_n13288_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X22 c1_n13188_n13100# m3_n7969_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X23 c1_n13188_n13100# m3_n2650_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X24 c1_n13188_n13100# m3_2669_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
C0 m3_2669_n13200# m3_2669_n7900# 3.28fF
C1 m3_7988_8000# m3_2669_8000# 2.73fF
C2 c1_n13188_n13100# m3_7988_n7900# 61.01fF
C3 m3_n7969_n13200# c1_n13188_n13100# 58.61fF
C4 c1_n13188_n13100# m3_n13288_n13200# 58.36fF
C5 m3_n7969_n13200# m3_n2650_n13200# 2.73fF
C6 c1_n13188_n13100# m3_n2650_2700# 58.86fF
C7 m3_n7969_n7900# m3_n13288_n7900# 2.73fF
C8 c1_n13188_n13100# m3_n7969_8000# 58.61fF
C9 m3_2669_2700# m3_n2650_2700# 2.73fF
C10 m3_2669_n2600# c1_n13188_n13100# 58.86fF
C11 m3_7988_n13200# m3_7988_n7900# 3.39fF
C12 c1_n13188_n13100# m3_n2650_n13200# 58.61fF
C13 m3_2669_2700# c1_n13188_n13100# 58.86fF
C14 m3_n2650_2700# m3_n7969_2700# 2.73fF
C15 c1_n13188_n13100# m3_n13288_n2600# 58.61fF
C16 c1_n13188_n13100# m3_n2650_n7900# 58.86fF
C17 c1_n13188_n13100# m3_n7969_2700# 58.86fF
C18 m3_2669_2700# m3_2669_n2600# 3.28fF
C19 m3_n2650_n2600# m3_n7969_n2600# 2.73fF
C20 m3_n7969_8000# m3_n7969_2700# 3.28fF
C21 m3_7988_n13200# c1_n13188_n13100# 60.75fF
C22 m3_n2650_n7900# m3_n2650_n13200# 3.28fF
C23 m3_n7969_n7900# m3_n7969_n2600# 3.28fF
C24 m3_n2650_8000# m3_n2650_2700# 3.28fF
C25 m3_7988_n2600# m3_7988_n7900# 3.39fF
C26 c1_n13188_n13100# m3_n2650_8000# 58.61fF
C27 m3_2669_n13200# c1_n13188_n13100# 58.61fF
C28 m3_n2650_8000# m3_n7969_8000# 2.73fF
C29 m3_7988_2700# c1_n13188_n13100# 61.01fF
C30 c1_n13188_n13100# m3_n13288_8000# 58.36fF
C31 m3_n13288_n7900# m3_n13288_n13200# 3.28fF
C32 c1_n13188_n13100# m3_7988_8000# 60.75fF
C33 m3_n13288_8000# m3_n7969_8000# 2.73fF
C34 m3_2669_n13200# m3_n2650_n13200# 2.73fF
C35 m3_2669_n7900# m3_7988_n7900# 2.73fF
C36 m3_2669_2700# m3_7988_2700# 2.73fF
C37 m3_7988_n2600# c1_n13188_n13100# 61.01fF
C38 c1_n13188_n13100# m3_n13288_n7900# 58.61fF
C39 c1_n13188_n13100# m3_n13288_2700# 58.61fF
C40 m3_7988_n2600# m3_2669_n2600# 2.73fF
C41 m3_n7969_n13200# m3_n7969_n7900# 3.28fF
C42 m3_7988_n13200# m3_2669_n13200# 2.73fF
C43 c1_n13188_n13100# m3_2669_8000# 58.61fF
C44 m3_n13288_n7900# m3_n13288_n2600# 3.28fF
C45 m3_n2650_n2600# m3_n2650_2700# 3.28fF
C46 c1_n13188_n13100# m3_2669_n7900# 58.86fF
C47 m3_n13288_2700# m3_n13288_n2600# 3.28fF
C48 m3_n13288_2700# m3_n7969_2700# 2.73fF
C49 c1_n13188_n13100# m3_n2650_n2600# 58.86fF
C50 m3_2669_n2600# m3_2669_n7900# 3.28fF
C51 c1_n13188_n13100# m3_n7969_n2600# 58.86fF
C52 m3_2669_2700# m3_2669_8000# 3.28fF
C53 m3_2669_n2600# m3_n2650_n2600# 2.73fF
C54 c1_n13188_n13100# m3_n7969_n7900# 58.86fF
C55 m3_7988_2700# m3_7988_8000# 3.39fF
C56 m3_n2650_n7900# m3_2669_n7900# 2.73fF
C57 m3_n2650_n7900# m3_n2650_n2600# 3.28fF
C58 m3_n13288_n2600# m3_n7969_n2600# 2.73fF
C59 m3_7988_2700# m3_7988_n2600# 3.39fF
C60 m3_n7969_n2600# m3_n7969_2700# 3.28fF
C61 m3_n13288_8000# m3_n13288_2700# 3.28fF
C62 m3_n2650_n7900# m3_n7969_n7900# 2.73fF
C63 m3_n7969_n13200# m3_n13288_n13200# 2.73fF
C64 m3_n2650_8000# m3_2669_8000# 2.73fF
C65 c1_n13188_n13100# VSUBS 2.51fF
C66 m3_7988_n13200# VSUBS 12.57fF
C67 m3_2669_n13200# VSUBS 12.37fF
C68 m3_n2650_n13200# VSUBS 12.37fF
C69 m3_n7969_n13200# VSUBS 12.37fF
C70 m3_n13288_n13200# VSUBS 12.37fF
C71 m3_7988_n7900# VSUBS 12.57fF
C72 m3_2669_n7900# VSUBS 12.37fF
C73 m3_n2650_n7900# VSUBS 12.37fF
C74 m3_n7969_n7900# VSUBS 12.37fF
C75 m3_n13288_n7900# VSUBS 12.37fF
C76 m3_7988_n2600# VSUBS 12.57fF
C77 m3_2669_n2600# VSUBS 12.37fF
C78 m3_n2650_n2600# VSUBS 12.37fF
C79 m3_n7969_n2600# VSUBS 12.37fF
C80 m3_n13288_n2600# VSUBS 12.37fF
C81 m3_7988_2700# VSUBS 12.57fF
C82 m3_2669_2700# VSUBS 12.37fF
C83 m3_n2650_2700# VSUBS 12.37fF
C84 m3_n7969_2700# VSUBS 12.37fF
C85 m3_n13288_2700# VSUBS 12.37fF
C86 m3_7988_8000# VSUBS 12.57fF
C87 m3_2669_8000# VSUBS 12.37fF
C88 m3_n2650_8000# VSUBS 12.37fF
C89 m3_n7969_8000# VSUBS 12.37fF
C90 m3_n13288_8000# VSUBS 12.37fF
.ends

.subckt cap1_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_MACBVW_0 VSUBS out out out out out out out out out out
+ out out out out out out out out out out out in out out out out sky130_fd_pr__cap_mim_m3_1_MACBVW
C0 in out 2.17fF
C1 in VSUBS -10.03fF
C2 out VSUBS 62.40fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WHJTNJ VSUBS m3_n4309_50# m3_n4309_n4250# c1_n4209_n4150#
+ c1_110_n4150# m3_10_n4250#
X0 c1_n4209_n4150# m3_n4309_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 c1_110_n4150# m3_10_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2 c1_n4209_n4150# m3_n4309_50# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 c1_110_n4150# m3_10_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
C0 m3_n4309_n4250# m3_n4309_50# 2.63fF
C1 m3_n4309_50# m3_10_n4250# 1.75fF
C2 c1_n4209_n4150# m3_n4309_50# 38.10fF
C3 c1_110_n4150# m3_10_n4250# 81.11fF
C4 c1_110_n4150# c1_n4209_n4150# 1.32fF
C5 m3_n4309_n4250# m3_10_n4250# 1.75fF
C6 m3_n4309_n4250# c1_n4209_n4150# 38.10fF
C7 c1_110_n4150# VSUBS 0.12fF
C8 c1_n4209_n4150# VSUBS 0.12fF
C9 m3_n4309_n4250# VSUBS 8.68fF
C10 m3_10_n4250# VSUBS 17.92fF
C11 m3_n4309_50# VSUBS 8.68fF
.ends

.subckt cap3_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_WHJTNJ_0 VSUBS out out in in out sky130_fd_pr__cap_mim_m3_1_WHJTNJ
C0 out in 3.21fF
C1 in VSUBS -8.91fF
C2 out VSUBS 3.92fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_W3JTNJ VSUBS m3_n6469_n2100# c1_n6369_n6300# m3_2169_n6400#
+ m3_n2150_n6400# c1_2269_n6300# m3_n6469_2200# m3_n2150_n2100# c1_n2050_n6300# m3_n2150_2200#
+ m3_n6469_n6400#
X0 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2 c1_n2050_n6300# m3_n2150_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 c1_n6369_n6300# m3_n6469_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X4 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X5 c1_n6369_n6300# m3_n6469_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X6 c1_n2050_n6300# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X7 c1_n2050_n6300# m3_n2150_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X8 c1_n6369_n6300# m3_n6469_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
C0 c1_n2050_n6300# m3_n2150_2200# 38.10fF
C1 m3_n6469_n2100# c1_n6369_n6300# 38.10fF
C2 m3_n6469_n6400# c1_n6369_n6300# 38.10fF
C3 m3_n6469_n2100# m3_n2150_n2100# 1.75fF
C4 m3_n2150_n2100# m3_n2150_n6400# 2.63fF
C5 m3_n6469_n2100# m3_n6469_2200# 2.63fF
C6 m3_2169_n6400# m3_n2150_n6400# 1.75fF
C7 m3_n2150_n2100# m3_n2150_2200# 2.63fF
C8 m3_n2150_2200# m3_n6469_2200# 1.75fF
C9 m3_2169_n6400# m3_n2150_2200# 1.75fF
C10 c1_2269_n6300# c1_n2050_n6300# 1.99fF
C11 c1_n6369_n6300# c1_n2050_n6300# 1.99fF
C12 m3_n2150_n2100# c1_n2050_n6300# 38.10fF
C13 c1_2269_n6300# m3_2169_n6400# 121.67fF
C14 c1_n6369_n6300# m3_n6469_2200# 38.10fF
C15 m3_2169_n6400# m3_n2150_n2100# 1.75fF
C16 m3_n6469_n6400# m3_n6469_n2100# 2.63fF
C17 m3_n6469_n6400# m3_n2150_n6400# 1.75fF
C18 m3_n2150_n6400# c1_n2050_n6300# 38.10fF
C19 c1_2269_n6300# VSUBS 0.16fF
C20 c1_n2050_n6300# VSUBS 0.16fF
C21 c1_n6369_n6300# VSUBS 0.16fF
C22 m3_n2150_n6400# VSUBS 8.68fF
C23 m3_n6469_n6400# VSUBS 8.68fF
C24 m3_n2150_n2100# VSUBS 8.68fF
C25 m3_n6469_n2100# VSUBS 8.68fF
C26 m3_2169_n6400# VSUBS 26.86fF
C27 m3_n2150_2200# VSUBS 8.68fF
C28 m3_n6469_2200# VSUBS 8.68fF
.ends

.subckt cap2_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_W3JTNJ_0 VSUBS out in out out in out out in out out sky130_fd_pr__cap_mim_m3_1_W3JTNJ
C0 in out 8.08fF
C1 in VSUBS -16.59fF
C2 out VSUBS 13.00fF
.ends

.subckt sky130_fd_pr__nfet_01v8_U2JGXT w_n226_n510# a_n118_n388# a_n88_n300# a_30_n300#
X0 a_30_n300# a_n118_n388# a_n88_n300# w_n226_n510# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
C0 a_n88_n300# a_n118_n388# 0.11fF
C1 a_n88_n300# a_30_n300# 0.61fF
C2 a_30_n300# w_n226_n510# 0.40fF
C3 a_n88_n300# w_n226_n510# 0.40fF
C4 a_n118_n388# w_n226_n510# 0.28fF
.ends

.subckt sky130_fd_pr__res_high_po_5p73_X44RQA a_n573_2292# w_n739_n2890# a_n573_n2724#
X0 a_n573_n2724# a_n573_2292# w_n739_n2890# sky130_fd_pr__res_high_po_5p73 l=2.292e+07u
C0 a_n573_n2724# w_n739_n2890# 1.98fF
C1 a_n573_2292# w_n739_n2890# 1.98fF
.ends

.subckt res_loop_filter vss out in
Xsky130_fd_pr__res_high_po_5p73_X44RQA_0 in vss out sky130_fd_pr__res_high_po_5p73_X44RQA
C0 out vss 3.87fF
C1 in vss 3.02fF
.ends

.subckt loop_filter_v2 vc_pex D0_cap in vss
Xcap1_loop_filter_0 vss vc_pex vss cap1_loop_filter
Xcap3_loop_filter_0 vss cap3_loop_filter_0/in vss cap3_loop_filter
Xcap2_loop_filter_0 vss in vss cap2_loop_filter
Xsky130_fd_pr__nfet_01v8_U2JGXT_0 vss D0_cap in cap3_loop_filter_0/in sky130_fd_pr__nfet_01v8_U2JGXT
Xres_loop_filter_0 vss res_loop_filter_2/out in res_loop_filter
Xres_loop_filter_1 vss res_loop_filter_2/out vc_pex res_loop_filter
Xres_loop_filter_2 vss res_loop_filter_2/out vc_pex res_loop_filter
C0 D0_cap in 0.07fF
C1 cap3_loop_filter_0/in in 0.79fF
C2 vc_pex in 0.18fF
C3 vc_pex vss -38.13fF
C4 res_loop_filter_2/out vss 8.49fF
C5 D0_cap vss 0.04fF
C6 in vss -18.54fF
C7 cap3_loop_filter_0/in vss -3.74fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4798MH VSUBS w_n311_n338# a_81_n156# a_111_n125# a_15_n125#
+ a_n173_n125# a_n111_n156# a_n15_n156# a_n81_n125#
X0 a_n81_n125# a_n111_n156# a_n173_n125# w_n311_n338# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n15_n156# a_n81_n125# w_n311_n338# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_81_n156# a_15_n125# w_n311_n338# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_111_n125# a_n173_n125# 0.08fF
C1 a_n15_n156# a_n111_n156# 0.02fF
C2 a_n15_n156# a_81_n156# 0.02fF
C3 a_n81_n125# a_15_n125# 0.36fF
C4 a_n81_n125# a_n173_n125# 0.36fF
C5 a_n173_n125# a_15_n125# 0.13fF
C6 a_111_n125# a_n81_n125# 0.13fF
C7 a_111_n125# a_15_n125# 0.36fF
C8 a_111_n125# VSUBS 0.03fF
C9 a_15_n125# VSUBS 0.03fF
C10 a_n81_n125# VSUBS 0.03fF
C11 a_n173_n125# VSUBS 0.03fF
C12 a_81_n156# VSUBS 0.05fF
C13 a_n15_n156# VSUBS 0.05fF
C14 a_n111_n156# VSUBS 0.05fF
C15 w_n311_n338# VSUBS 1.56fF
.ends

.subckt sky130_fd_pr__nfet_01v8_BHR94T a_n15_n151# w_n311_n335# a_81_n151# a_111_n125#
+ a_15_n125# a_n173_n125# a_n111_n151# a_n81_n125#
X0 a_111_n125# a_81_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n15_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_81_n151# a_n15_n151# 0.02fF
C1 a_15_n125# a_111_n125# 0.36fF
C2 a_n15_n151# a_n111_n151# 0.02fF
C3 a_15_n125# a_n173_n125# 0.13fF
C4 a_n173_n125# a_111_n125# 0.08fF
C5 a_15_n125# a_n81_n125# 0.36fF
C6 a_n81_n125# a_111_n125# 0.13fF
C7 a_n81_n125# a_n173_n125# 0.36fF
C8 a_111_n125# w_n311_n335# 0.04fF
C9 a_15_n125# w_n311_n335# 0.04fF
C10 a_n81_n125# w_n311_n335# 0.04fF
C11 a_n173_n125# w_n311_n335# 0.04fF
C12 a_81_n151# w_n311_n335# 0.05fF
C13 a_n15_n151# w_n311_n335# 0.05fF
C14 a_n111_n151# w_n311_n335# 0.05fF
.ends

.subckt trans_gate m1_187_n605# vss m1_45_n513# vdd
Xsky130_fd_pr__pfet_01v8_4798MH_0 vss vdd vss m1_187_n605# m1_45_n513# m1_45_n513#
+ vss vss m1_187_n605# sky130_fd_pr__pfet_01v8_4798MH
Xsky130_fd_pr__nfet_01v8_BHR94T_0 vdd vss vdd m1_187_n605# m1_45_n513# m1_45_n513#
+ vdd m1_187_n605# sky130_fd_pr__nfet_01v8_BHR94T
C0 m1_187_n605# m1_45_n513# 0.36fF
C1 vdd m1_45_n513# 0.69fF
C2 vdd m1_187_n605# 0.55fF
C3 m1_187_n605# vss 0.73fF
C4 m1_45_n513# vss 1.10fF
C5 vdd vss 2.55fF
.ends

.subckt sky130_fd_pr__pfet_01v8_7KT7MH VSUBS a_n111_n186# a_111_n125# a_15_n125# a_n173_n125#
+ w_n311_n344# a_n81_n125#
X0 a_n81_n125# a_n111_n186# a_n173_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n111_n186# a_n81_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_n111_n186# a_15_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n173_n125# w_n311_n344# 0.14fF
C1 w_n311_n344# a_111_n125# 0.14fF
C2 a_n81_n125# a_15_n125# 0.36fF
C3 a_n173_n125# a_15_n125# 0.13fF
C4 a_111_n125# a_15_n125# 0.36fF
C5 a_n173_n125# a_n81_n125# 0.36fF
C6 w_n311_n344# a_15_n125# 0.09fF
C7 a_111_n125# a_n81_n125# 0.13fF
C8 a_n173_n125# a_111_n125# 0.08fF
C9 w_n311_n344# a_n81_n125# 0.09fF
C10 a_111_n125# VSUBS 0.03fF
C11 a_15_n125# VSUBS 0.03fF
C12 a_n81_n125# VSUBS 0.03fF
C13 a_n173_n125# VSUBS 0.03fF
C14 a_n111_n186# VSUBS 0.26fF
C15 w_n311_n344# VSUBS 2.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS6QM w_n311_n335# a_111_n125# a_15_n125# a_n173_n125#
+ a_n111_n151# a_n81_n125#
X0 a_111_n125# a_n111_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n111_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_15_n125# a_111_n125# 0.36fF
C1 a_n81_n125# a_111_n125# 0.13fF
C2 a_n173_n125# a_111_n125# 0.08fF
C3 a_n81_n125# a_15_n125# 0.36fF
C4 a_n173_n125# a_15_n125# 0.13fF
C5 a_n81_n125# a_n173_n125# 0.36fF
C6 a_111_n125# w_n311_n335# 0.17fF
C7 a_15_n125# w_n311_n335# 0.12fF
C8 a_n81_n125# w_n311_n335# 0.12fF
C9 a_n173_n125# w_n311_n335# 0.17fF
C10 a_n111_n151# w_n311_n335# 0.25fF
.ends

.subckt inverter_cp_x1 out in vss vdd
Xsky130_fd_pr__pfet_01v8_7KT7MH_0 vss in out vdd vdd vdd out sky130_fd_pr__pfet_01v8_7KT7MH
Xsky130_fd_pr__nfet_01v8_2BS6QM_0 vss out vss vss in out sky130_fd_pr__nfet_01v8_2BS6QM
C0 out in 0.32fF
C1 vdd out 0.10fF
C2 out vss 0.77fF
C3 in vss 0.95fF
C4 vdd vss 3.13fF
.ends

.subckt clock_inverter vss inverter_cp_x1_2/in CLK vdd inverter_cp_x1_0/out CLK_d
+ nCLK_d
Xtrans_gate_0 nCLK_d vss inverter_cp_x1_0/out vdd trans_gate
Xinverter_cp_x1_0 inverter_cp_x1_0/out CLK vss vdd inverter_cp_x1
Xinverter_cp_x1_1 inverter_cp_x1_2/in CLK vss vdd inverter_cp_x1
Xinverter_cp_x1_2 CLK_d inverter_cp_x1_2/in vss vdd inverter_cp_x1
C0 CLK_d inverter_cp_x1_2/in 0.12fF
C1 CLK_d vdd 0.03fF
C2 inverter_cp_x1_0/out vdd 0.21fF
C3 inverter_cp_x1_2/in vdd 0.21fF
C4 inverter_cp_x1_0/out nCLK_d 0.11fF
C5 vdd nCLK_d 0.03fF
C6 inverter_cp_x1_0/out CLK 0.31fF
C7 inverter_cp_x1_2/in CLK 0.31fF
C8 vdd CLK 0.36fF
C9 CLK_d vss 0.96fF
C10 inverter_cp_x1_2/in vss 2.01fF
C11 inverter_cp_x1_0/out vss 1.69fF
C12 CLK vss 3.03fF
C13 vdd vss 15.46fF
C14 nCLK_d vss 1.23fF
.ends

.subckt sky130_fd_pr__pfet_01v8_MJG8BZ VSUBS a_n125_n95# a_63_n95# w_n263_n314# a_n33_n95#
+ a_n63_n192#
X0 a_63_n95# a_n63_n192# a_n33_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n33_n95# a_n63_n192# a_n125_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
C0 w_n263_n314# a_63_n95# 0.11fF
C1 w_n263_n314# a_n125_n95# 0.11fF
C2 a_63_n95# a_n125_n95# 0.10fF
C3 w_n263_n314# a_n33_n95# 0.08fF
C4 a_n33_n95# a_63_n95# 0.28fF
C5 a_n33_n95# a_n125_n95# 0.28fF
C6 a_63_n95# VSUBS 0.03fF
C7 a_n33_n95# VSUBS 0.03fF
C8 a_n125_n95# VSUBS 0.03fF
C9 a_n63_n192# VSUBS 0.20fF
C10 w_n263_n314# VSUBS 1.80fF
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS854 w_n311_n335# a_n129_n213# a_111_n125# a_15_n125#
+ a_n173_n125# a_n81_n125#
X0 a_111_n125# a_n129_n213# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n129_n213# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n129_n213# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_15_n125# a_n173_n125# 0.13fF
C1 a_n129_n213# a_111_n125# 0.01fF
C2 a_n129_n213# a_n81_n125# 0.10fF
C3 a_111_n125# a_n81_n125# 0.13fF
C4 a_n129_n213# a_15_n125# 0.10fF
C5 a_15_n125# a_111_n125# 0.36fF
C6 a_15_n125# a_n81_n125# 0.36fF
C7 a_n129_n213# a_n173_n125# 0.02fF
C8 a_111_n125# a_n173_n125# 0.08fF
C9 a_n173_n125# a_n81_n125# 0.36fF
C10 a_111_n125# w_n311_n335# 0.05fF
C11 a_15_n125# w_n311_n335# 0.05fF
C12 a_n81_n125# w_n311_n335# 0.05fF
C13 a_n173_n125# w_n311_n335# 0.05fF
C14 a_n129_n213# w_n311_n335# 0.49fF
.ends

.subckt sky130_fd_pr__nfet_01v8_KU9PSX a_n125_n95# a_n33_n95# a_n81_n183# w_n263_n305#
X0 a_n33_n95# a_n81_n183# a_n125_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n125_n95# a_n81_n183# a_n33_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
C0 a_n81_n183# a_n33_n95# 0.10fF
C1 a_n81_n183# a_n125_n95# 0.16fF
C2 a_n125_n95# a_n33_n95# 0.88fF
C3 a_n33_n95# w_n263_n305# 0.07fF
C4 a_n125_n95# w_n263_n305# 0.13fF
C5 a_n81_n183# w_n263_n305# 0.31fF
.ends

.subckt latch_diff m1_657_280# nQ Q vss CLK vdd nD D
Xsky130_fd_pr__pfet_01v8_MJG8BZ_0 vss vdd vdd vdd nQ Q sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__pfet_01v8_MJG8BZ_1 vss vdd vdd vdd Q nQ sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__nfet_01v8_2BS854_0 vss CLK vss m1_657_280# m1_657_280# vss sky130_fd_pr__nfet_01v8_2BS854
Xsky130_fd_pr__nfet_01v8_KU9PSX_0 m1_657_280# Q nD vss sky130_fd_pr__nfet_01v8_KU9PSX
Xsky130_fd_pr__nfet_01v8_KU9PSX_1 m1_657_280# nQ D vss sky130_fd_pr__nfet_01v8_KU9PSX
C0 Q nQ 0.93fF
C1 nD Q 0.05fF
C2 nD nQ 0.05fF
C3 vdd Q 0.16fF
C4 vdd nQ 0.16fF
C5 D Q 0.05fF
C6 m1_657_280# Q 0.94fF
C7 D nQ 0.05fF
C8 m1_657_280# CLK 0.24fF
C9 m1_657_280# nQ 1.41fF
C10 D vss 0.53fF
C11 m1_657_280# vss 1.88fF
C12 nD vss 0.16fF
C13 CLK vss 0.87fF
C14 Q vss -0.55fF
C15 nQ vss 1.16fF
C16 vdd vss 5.98fF
.ends

.subckt DFlipFlop latch_diff_0/m1_657_280# vdd vss latch_diff_1/D clock_inverter_0/inverter_cp_x1_2/in
+ nQ nCLK latch_diff_0/nD Q latch_diff_1/nD D latch_diff_1/m1_657_280# latch_diff_0/D
+ CLK clock_inverter_0/inverter_cp_x1_0/out
Xclock_inverter_0 vss clock_inverter_0/inverter_cp_x1_2/in D vdd clock_inverter_0/inverter_cp_x1_0/out
+ latch_diff_0/D latch_diff_0/nD clock_inverter
Xlatch_diff_0 latch_diff_0/m1_657_280# latch_diff_1/nD latch_diff_1/D vss CLK vdd
+ latch_diff_0/nD latch_diff_0/D latch_diff
Xlatch_diff_1 latch_diff_1/m1_657_280# nQ Q vss nCLK vdd latch_diff_1/nD latch_diff_1/D
+ latch_diff
C0 latch_diff_1/D latch_diff_1/nD 0.33fF
C1 latch_diff_1/D latch_diff_0/D 0.11fF
C2 vdd latch_diff_1/nD 0.02fF
C3 vdd latch_diff_0/D 0.09fF
C4 latch_diff_1/m1_657_280# latch_diff_0/m1_657_280# 0.18fF
C5 latch_diff_1/m1_657_280# latch_diff_1/nD 0.42fF
C6 latch_diff_0/m1_657_280# latch_diff_1/nD 0.14fF
C7 latch_diff_0/m1_657_280# latch_diff_0/D 0.37fF
C8 latch_diff_0/D latch_diff_1/nD 0.04fF
C9 latch_diff_1/D latch_diff_0/nD 0.41fF
C10 clock_inverter_0/inverter_cp_x1_0/out vdd 0.03fF
C11 vdd latch_diff_0/nD 0.14fF
C12 nQ latch_diff_1/D 0.11fF
C13 Q latch_diff_1/nD 0.01fF
C14 latch_diff_1/D vdd 0.01fF
C15 latch_diff_0/m1_657_280# latch_diff_0/nD 0.38fF
C16 latch_diff_1/m1_657_280# latch_diff_1/D 0.32fF
C17 latch_diff_1/D latch_diff_0/m1_657_280# 0.43fF
C18 nQ latch_diff_1/nD 0.08fF
C19 latch_diff_1/m1_657_280# vss 0.64fF
C20 nCLK vss 0.83fF
C21 Q vss -0.92fF
C22 nQ vss 0.57fF
C23 latch_diff_0/m1_657_280# vss 0.69fF
C24 CLK vss 0.83fF
C25 latch_diff_1/D vss -0.33fF
C26 latch_diff_1/nD vss 1.83fF
C27 latch_diff_0/D vss 1.29fF
C28 clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C29 clock_inverter_0/inverter_cp_x1_0/out vss 1.63fF
C30 D vss 3.27fF
C31 vdd vss 31.85fF
C32 latch_diff_0/nD vss 1.53fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ZP3U9B VSUBS a_n221_n84# a_159_n84# w_n359_n303# a_n63_n110#
+ a_n129_n84# a_33_n110# a_n159_n110# a_63_n84# a_129_n110# a_n33_n84#
X0 a_n129_n84# a_n159_n110# a_n221_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_63_n84# a_33_n110# a_n33_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_n33_n84# a_n63_n110# a_n129_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_159_n84# a_129_n110# a_63_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_n221_n84# w_n359_n303# 0.08fF
C1 a_159_n84# a_n221_n84# 0.04fF
C2 a_n221_n84# a_n33_n84# 0.09fF
C3 a_33_n110# a_129_n110# 0.02fF
C4 a_63_n84# w_n359_n303# 0.06fF
C5 a_63_n84# a_159_n84# 0.24fF
C6 a_63_n84# a_n33_n84# 0.24fF
C7 a_n63_n110# a_n159_n110# 0.02fF
C8 a_n129_n84# a_n221_n84# 0.24fF
C9 a_n129_n84# a_63_n84# 0.09fF
C10 a_159_n84# w_n359_n303# 0.08fF
C11 w_n359_n303# a_n33_n84# 0.05fF
C12 a_159_n84# a_n33_n84# 0.09fF
C13 a_n129_n84# w_n359_n303# 0.06fF
C14 a_n63_n110# a_33_n110# 0.02fF
C15 a_n129_n84# a_159_n84# 0.05fF
C16 a_n129_n84# a_n33_n84# 0.24fF
C17 a_63_n84# a_n221_n84# 0.05fF
C18 a_159_n84# VSUBS 0.03fF
C19 a_63_n84# VSUBS 0.03fF
C20 a_n33_n84# VSUBS 0.03fF
C21 a_n129_n84# VSUBS 0.03fF
C22 a_n221_n84# VSUBS 0.03fF
C23 a_129_n110# VSUBS 0.05fF
C24 a_33_n110# VSUBS 0.05fF
C25 a_n63_n110# VSUBS 0.05fF
C26 a_n159_n110# VSUBS 0.05fF
C27 w_n359_n303# VSUBS 2.19fF
.ends

.subckt sky130_fd_pr__nfet_01v8_DXA56D w_n359_n252# a_n33_n42# a_129_n68# a_n159_n68#
+ a_n221_n42# a_159_n42# a_n129_n42# a_33_n68# a_n63_n68# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n129_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_159_n42# a_129_n68# a_63_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_n129_n42# a_n159_n68# a_n221_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n159_n68# a_n63_n68# 0.02fF
C1 a_n33_n42# a_63_n42# 0.12fF
C2 a_159_n42# a_n129_n42# 0.03fF
C3 a_n129_n42# a_n221_n42# 0.12fF
C4 a_159_n42# a_n221_n42# 0.02fF
C5 a_33_n68# a_129_n68# 0.02fF
C6 a_n63_n68# a_33_n68# 0.02fF
C7 a_n129_n42# a_63_n42# 0.05fF
C8 a_n129_n42# a_n33_n42# 0.12fF
C9 a_159_n42# a_63_n42# 0.12fF
C10 a_159_n42# a_n33_n42# 0.05fF
C11 a_n221_n42# a_63_n42# 0.03fF
C12 a_n33_n42# a_n221_n42# 0.05fF
C13 a_159_n42# w_n359_n252# 0.07fF
C14 a_63_n42# w_n359_n252# 0.06fF
C15 a_n33_n42# w_n359_n252# 0.06fF
C16 a_n129_n42# w_n359_n252# 0.06fF
C17 a_n221_n42# w_n359_n252# 0.07fF
C18 a_129_n68# w_n359_n252# 0.05fF
C19 a_33_n68# w_n359_n252# 0.05fF
C20 a_n63_n68# w_n359_n252# 0.05fF
C21 a_n159_n68# w_n359_n252# 0.05fF
.ends

.subckt inverter_min_x4 in vss out vdd
Xsky130_fd_pr__pfet_01v8_ZP3U9B_0 vss out out vdd in vdd in in vdd in out sky130_fd_pr__pfet_01v8_ZP3U9B
Xsky130_fd_pr__nfet_01v8_DXA56D_0 vss out in in out out vss in in vss sky130_fd_pr__nfet_01v8_DXA56D
C0 vdd out 0.62fF
C1 in out 0.67fF
C2 vdd in 0.33fF
C3 out vss 0.66fF
C4 in vss 1.89fF
C5 vdd vss 3.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_5RJ8EK a_n33_n42# a_33_n68# w_n263_n252# a_n63_n68#
+ a_n125_n42# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n125_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_63_n42# a_n125_n42# 0.05fF
C1 a_n33_n42# a_n125_n42# 0.12fF
C2 a_n33_n42# a_63_n42# 0.12fF
C3 a_33_n68# a_n63_n68# 0.02fF
C4 a_63_n42# w_n263_n252# 0.09fF
C5 a_n33_n42# w_n263_n252# 0.07fF
C6 a_n125_n42# w_n263_n252# 0.09fF
C7 a_33_n68# w_n263_n252# 0.05fF
C8 a_n63_n68# w_n263_n252# 0.05fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ZPB9BB VSUBS a_n63_n110# a_33_n110# a_n125_n84# a_63_n84#
+ w_n263_n303# a_n33_n84#
X0 a_63_n84# a_33_n110# a_n33_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_n33_n84# a_n63_n110# a_n125_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_63_n84# w_n263_n303# 0.10fF
C1 a_63_n84# a_n33_n84# 0.24fF
C2 a_n33_n84# w_n263_n303# 0.07fF
C3 a_63_n84# a_n125_n84# 0.09fF
C4 a_n125_n84# w_n263_n303# 0.10fF
C5 a_n63_n110# a_33_n110# 0.02fF
C6 a_n125_n84# a_n33_n84# 0.24fF
C7 a_63_n84# VSUBS 0.03fF
C8 a_n33_n84# VSUBS 0.03fF
C9 a_n125_n84# VSUBS 0.03fF
C10 a_33_n110# VSUBS 0.05fF
C11 a_n63_n110# VSUBS 0.05fF
C12 w_n263_n303# VSUBS 1.74fF
.ends

.subckt inverter_min_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_5RJ8EK_0 vss in vss in out out sky130_fd_pr__nfet_01v8_5RJ8EK
Xsky130_fd_pr__pfet_01v8_ZPB9BB_0 vss in in out out vdd vdd sky130_fd_pr__pfet_01v8_ZPB9BB
C0 vdd in 0.01fF
C1 out in 0.30fF
C2 vdd out 0.15fF
C3 vdd vss 2.93fF
C4 out vss 0.66fF
C5 in vss 0.72fF
.ends

.subckt div_by_2 vdd vss nout_div CLK_2 nCLK_2 o1 o2 CLK out_div
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vdd vss DFlipFlop_0/latch_diff_1/D
+ DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in nout_div DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_0/nD
+ out_div DFlipFlop_0/latch_diff_1/nD nout_div DFlipFlop_0/latch_diff_1/m1_657_280#
+ DFlipFlop_0/latch_diff_0/D DFlipFlop_0/CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
Xclock_inverter_0 vss clock_inverter_0/inverter_cp_x1_2/in CLK vdd clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_0/CLK DFlipFlop_0/nCLK clock_inverter
Xinverter_min_x4_1 o2 vss nCLK_2 vdd inverter_min_x4
Xinverter_min_x4_0 o1 vss CLK_2 vdd inverter_min_x4
Xinverter_min_x2_0 nout_div o2 vss vdd inverter_min_x2
Xinverter_min_x2_1 out_div o1 vss vdd inverter_min_x2
C0 o2 vdd 0.14fF
C1 nout_div DFlipFlop_0/latch_diff_0/D 0.09fF
C2 DFlipFlop_0/latch_diff_1/m1_657_280# DFlipFlop_0/nCLK 0.26fF
C3 nout_div DFlipFlop_0/latch_diff_1/D 0.64fF
C4 vdd DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C5 o1 vdd 0.14fF
C6 nCLK_2 vdd 0.08fF
C7 o2 DFlipFlop_0/latch_diff_1/m1_657_280# 0.02fF
C8 vdd nout_div 0.16fF
C9 o1 CLK_2 0.11fF
C10 DFlipFlop_0/latch_diff_1/nD nout_div 1.18fF
C11 DFlipFlop_0/latch_diff_0/nD nout_div 0.07fF
C12 DFlipFlop_0/CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.29fF
C13 DFlipFlop_0/CLK DFlipFlop_0/latch_diff_1/D -0.48fF
C14 vdd CLK_2 0.08fF
C15 nout_div DFlipFlop_0/CLK 0.42fF
C16 vdd DFlipFlop_0/CLK 0.40fF
C17 DFlipFlop_0/latch_diff_1/m1_657_280# o1 0.02fF
C18 nout_div DFlipFlop_0/latch_diff_0/m1_657_280# 0.24fF
C19 DFlipFlop_0/latch_diff_0/D DFlipFlop_0/nCLK 0.13fF
C20 DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/CLK 0.11fF
C21 DFlipFlop_0/latch_diff_0/nD DFlipFlop_0/CLK 0.12fF
C22 clock_inverter_0/inverter_cp_x1_0/out vdd 0.10fF
C23 DFlipFlop_0/latch_diff_1/m1_657_280# nout_div 0.21fF
C24 out_div o1 0.01fF
C25 DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_1/D 0.08fF
C26 DFlipFlop_0/CLK DFlipFlop_0/latch_diff_0/m1_657_280# 0.26fF
C27 out_div nout_div 0.22fF
C28 out_div vdd 0.03fF
C29 nout_div DFlipFlop_0/nCLK 0.43fF
C30 vdd DFlipFlop_0/nCLK 0.30fF
C31 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_0/nCLK 0.46fF
C32 DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/nCLK -0.09fF
C33 nCLK_2 o2 0.11fF
C34 CLK_2 vss 1.08fF
C35 o1 vss 2.21fF
C36 nCLK_2 vss 1.08fF
C37 o2 vss 2.21fF
C38 DFlipFlop_0/CLK vss 1.03fF
C39 clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C40 clock_inverter_0/inverter_cp_x1_0/out vss 1.64fF
C41 CLK vss 3.27fF
C42 DFlipFlop_0/nCLK vss 1.55fF
C43 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.63fF
C44 out_div vss -0.77fF
C45 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C46 DFlipFlop_0/latch_diff_1/D vss -1.72fF
C47 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C48 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C49 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C50 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.59fF
C51 nout_div vss 4.41fF
C52 vdd vss 62.89fF
C53 DFlipFlop_0/latch_diff_0/nD vss 0.94fF
.ends

.subckt trans_gate_mux2to8 in vss out en_pos en_neg vdd
Xsky130_fd_pr__pfet_01v8_4798MH_0 vss vdd en_neg in out out en_neg en_neg in sky130_fd_pr__pfet_01v8_4798MH
Xsky130_fd_pr__nfet_01v8_BHR94T_0 en_pos vss en_pos in out out en_pos in sky130_fd_pr__nfet_01v8_BHR94T
C0 en_neg in 0.28fF
C1 out en_neg 0.07fF
C2 en_neg en_pos 0.04fF
C3 out in 0.36fF
C4 in en_pos 0.07fF
C5 vdd in 0.05fF
C6 out en_pos 0.27fF
C7 out vdd 0.27fF
C8 vdd vss 2.08fF
C9 in vss 1.12fF
C10 out vss 0.87fF
C11 en_pos vss 0.29fF
C12 en_neg vss 0.31fF
.ends

.subckt mux2to1 vss select_0_neg out_a_0 out_a_1 select_0 vdd in_a
Xtrans_gate_mux2to8_0 in_a vss out_a_0 select_0_neg select_0 vdd trans_gate_mux2to8
Xtrans_gate_mux2to8_1 in_a vss out_a_1 select_0 select_0_neg vdd trans_gate_mux2to8
C0 out_a_1 in_a 0.08fF
C1 select_0 select_0_neg 0.17fF
C2 vdd out_a_0 0.06fF
C3 out_a_0 select_0_neg 0.05fF
C4 in_a select_0 0.31fF
C5 vdd in_a 0.02fF
C6 in_a select_0_neg 0.11fF
C7 in_a out_a_0 0.08fF
C8 out_a_1 select_0 0.14fF
C9 vdd out_a_1 0.06fF
C10 out_a_1 vss 0.99fF
C11 vdd vss 4.78fF
C12 in_a vss 2.00fF
C13 out_a_0 vss 0.99fF
C14 select_0_neg vss 1.15fF
C15 select_0 vss 0.97fF
.ends

.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X a_194_125# a_355_368# a_455_87#
X0 X B a_455_87# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 X a_194_125# a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_194_125# B a_158_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_158_392# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_355_368# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_194_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 a_455_87# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND B a_194_125# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X9 VGND a_194_125# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
C0 a_194_125# B 0.57fF
C1 a_194_125# X 0.29fF
C2 a_194_125# VPWR 0.33fF
C3 A VGND 0.31fF
C4 a_158_392# a_194_125# 0.06fF
C5 a_194_125# a_355_368# 0.51fF
C6 B X 0.13fF
C7 B VPWR 0.09fF
C8 B a_355_368# 0.08fF
C9 X VPWR 0.07fF
C10 X a_355_368# 0.17fF
C11 VPWR a_355_368# 0.37fF
C12 A a_194_125# 0.18fF
C13 VPWR VPB 0.06fF
C14 A B 0.28fF
C15 VGND a_194_125# 0.25fF
C16 VGND B 0.10fF
C17 A VPWR 0.15fF
C18 A a_355_368# 0.02fF
C19 VGND X 0.28fF
C20 VGND VPWR 0.01fF
C21 VGND VNB 0.78fF
C22 X VNB 0.21fF
C23 VPWR VNB 0.78fF
C24 B VNB 0.56fF
C25 A VNB 0.70fF
C26 VPB VNB 0.77fF
C27 a_355_368# VNB 0.08fF
C28 a_194_125# VNB 0.40fF
.ends

.subckt sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X a_143_136# a_56_136#
X0 VGND B a_143_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 X a_56_136# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VPWR B a_56_136# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_143_136# A a_56_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_56_136# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 X a_56_136# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
C0 A VGND 0.21fF
C1 X VGND 0.15fF
C2 VPWR A 0.07fF
C3 VPWR X 0.20fF
C4 B a_56_136# 0.30fF
C5 B VGND 0.03fF
C6 B VPWR 0.02fF
C7 a_56_136# VGND 0.06fF
C8 B A 0.08fF
C9 VPWR a_56_136# 0.57fF
C10 B X 0.02fF
C11 A a_56_136# 0.17fF
C12 a_56_136# X 0.26fF
C13 VPB VPWR 0.04fF
C14 VGND VNB 0.50fF
C15 X VNB 0.23fF
C16 VPWR VNB 0.50fF
C17 B VNB 0.24fF
C18 A VNB 0.36fF
C19 VPB VNB 0.48fF
C20 a_56_136# VNB 0.38fF
.ends

.subckt sky130_fd_sc_hs__or2_1 A B VGND VNB VPB VPWR X a_152_368# a_63_368#
X0 VPWR A a_152_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_152_368# B a_63_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 X a_63_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 X a_63_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_63_368# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X5 VGND A a_63_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
C0 VGND B 0.11fF
C1 X VGND 0.16fF
C2 VPWR A 0.05fF
C3 VGND a_63_368# 0.27fF
C4 A B 0.10fF
C5 X A 0.02fF
C6 a_63_368# A 0.28fF
C7 VPWR B 0.01fF
C8 X VPWR 0.18fF
C9 VPB VPWR 0.04fF
C10 VPWR a_63_368# 0.29fF
C11 a_63_368# B 0.14fF
C12 X a_63_368# 0.33fF
C13 a_152_368# a_63_368# 0.03fF
C14 VGND VNB 0.53fF
C15 X VNB 0.24fF
C16 A VNB 0.21fF
C17 B VNB 0.31fF
C18 VPWR VNB 0.46fF
C19 VPB VNB 0.48fF
C20 a_63_368# VNB 0.37fF
.ends

.subckt div_by_5 nCLK DFlipFlop_0/latch_diff_1/nD DFlipFlop_2/latch_diff_0/nD vss
+ Q1 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in CLK DFlipFlop_0/Q vdd DFlipFlop_2/latch_diff_1/D
+ DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out sky130_fd_sc_hs__and2_1_0/a_56_136#
+ DFlipFlop_3/latch_diff_0/D DFlipFlop_3/latch_diff_1/nD DFlipFlop_1/latch_diff_1/nD
+ DFlipFlop_1/latch_diff_0/nD DFlipFlop_2/latch_diff_0/m1_657_280# CLK_5 Q1_shift
+ nQ2 DFlipFlop_0/latch_diff_0/D DFlipFlop_2/D DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_1/latch_diff_1/D DFlipFlop_1/D nQ0 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_2/latch_diff_1/nD Q0 DFlipFlop_0/D DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_0/latch_diff_1/D DFlipFlop_0/latch_diff_0/nD DFlipFlop_2/nQ DFlipFlop_2/latch_diff_0/D
+ DFlipFlop_3/latch_diff_1/D sky130_fd_sc_hs__or2_1_0/a_152_368# sky130_fd_sc_hs__and2_1_1/a_56_136#
+ DFlipFlop_3/nQ sky130_fd_sc_hs__and2_1_0/a_143_136#
Xsky130_fd_sc_hs__xor2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_2/D sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ sky130_fd_sc_hs__xor2_1_0/a_355_368# sky130_fd_sc_hs__xor2_1_0/a_455_87# sky130_fd_sc_hs__xor2_1
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vdd vss DFlipFlop_0/latch_diff_1/D
+ DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in nQ2 nCLK DFlipFlop_0/latch_diff_0/nD
+ DFlipFlop_0/Q DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/D DFlipFlop_0/latch_diff_1/m1_657_280#
+ DFlipFlop_0/latch_diff_0/D CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_2 DFlipFlop_2/latch_diff_0/m1_657_280# vdd vss DFlipFlop_2/latch_diff_1/D
+ DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_2/nQ nCLK DFlipFlop_2/latch_diff_0/nD
+ Q1 DFlipFlop_2/latch_diff_1/nD DFlipFlop_2/D DFlipFlop_2/latch_diff_1/m1_657_280#
+ DFlipFlop_2/latch_diff_0/D CLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_1 DFlipFlop_1/latch_diff_0/m1_657_280# vdd vss DFlipFlop_1/latch_diff_1/D
+ DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in nQ0 nCLK DFlipFlop_1/latch_diff_0/nD
+ Q0 DFlipFlop_1/latch_diff_1/nD DFlipFlop_1/D DFlipFlop_1/latch_diff_1/m1_657_280#
+ DFlipFlop_1/latch_diff_0/D CLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_3 DFlipFlop_3/latch_diff_0/m1_657_280# vdd vss DFlipFlop_3/latch_diff_1/D
+ DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_3/nQ CLK DFlipFlop_3/latch_diff_0/nD
+ Q1_shift DFlipFlop_3/latch_diff_1/nD Q1 DFlipFlop_3/latch_diff_1/m1_657_280# DFlipFlop_3/latch_diff_0/D
+ nCLK DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop
Xsky130_fd_sc_hs__and2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_0/D sky130_fd_sc_hs__and2_1_0/a_143_136#
+ sky130_fd_sc_hs__and2_1_0/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__and2_1_1 nQ2 nQ0 vss vss vdd vdd DFlipFlop_1/D sky130_fd_sc_hs__and2_1_1/a_143_136#
+ sky130_fd_sc_hs__and2_1_1/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__or2_1_0 Q1 Q1_shift vss vss vdd vdd CLK_5 sky130_fd_sc_hs__or2_1_0/a_152_368#
+ sky130_fd_sc_hs__or2_1_0/a_63_368# sky130_fd_sc_hs__or2_1
C0 sky130_fd_sc_hs__and2_1_1/a_56_136# vdd 0.04fF
C1 DFlipFlop_0/latch_diff_1/D Q0 0.23fF
C2 nQ0 nCLK 0.09fF
C3 Q1_shift vdd 0.10fF
C4 Q1 DFlipFlop_1/D 0.03fF
C5 Q0 DFlipFlop_1/D 0.07fF
C6 DFlipFlop_2/latch_diff_1/D Q1 0.23fF
C7 Q0 DFlipFlop_1/latch_diff_1/m1_657_280# 0.01fF
C8 Q1 DFlipFlop_1/latch_diff_1/nD 0.10fF
C9 DFlipFlop_1/latch_diff_1/nD Q0 0.21fF
C10 Q1 Q0 9.65fF
C11 DFlipFlop_2/D vdd 0.07fF
C12 CLK DFlipFlop_2/latch_diff_1/nD 0.09fF
C13 sky130_fd_sc_hs__or2_1_0/a_152_368# Q1_shift -0.04fF
C14 CLK DFlipFlop_3/latch_diff_1/D 0.08fF
C15 DFlipFlop_1/D nCLK 0.14fF
C16 DFlipFlop_2/latch_diff_1/D nCLK 0.08fF
C17 DFlipFlop_1/latch_diff_1/m1_657_280# nCLK 0.28fF
C18 DFlipFlop_1/latch_diff_1/nD nCLK 0.16fF
C19 Q1 nCLK -0.01fF
C20 Q0 nCLK 0.20fF
C21 DFlipFlop_0/latch_diff_0/m1_657_280# CLK 0.28fF
C22 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vdd 0.03fF
C23 DFlipFlop_3/nQ Q1_shift 0.04fF
C24 Q1 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in 0.21fF
C25 nQ0 vdd 0.11fF
C26 Q0 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in 0.42fF
C27 Q0 sky130_fd_sc_hs__xor2_1_0/a_355_368# 0.03fF
C28 Q1 DFlipFlop_0/D 0.13fF
C29 Q1 sky130_fd_sc_hs__and2_1_0/a_56_136# 0.14fF
C30 DFlipFlop_0/D Q0 0.39fF
C31 DFlipFlop_1/latch_diff_1/D CLK 0.14fF
C32 Q0 sky130_fd_sc_hs__and2_1_0/a_56_136# 0.17fF
C33 CLK DFlipFlop_2/latch_diff_0/m1_657_280# 0.28fF
C34 CLK DFlipFlop_1/latch_diff_0/nD 0.08fF
C35 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in nCLK 0.14fF
C36 DFlipFlop_0/latch_diff_1/m1_657_280# nQ2 0.05fF
C37 Q1 DFlipFlop_0/Q 0.13fF
C38 Q0 DFlipFlop_0/Q 0.21fF
C39 DFlipFlop_1/D vdd 0.25fF
C40 DFlipFlop_3/latch_diff_1/nD CLK 0.16fF
C41 DFlipFlop_3/latch_diff_1/m1_657_280# CLK 0.27fF
C42 DFlipFlop_2/D sky130_fd_sc_hs__xor2_1_0/a_194_125# 0.08fF
C43 Q1 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out 0.15fF
C44 Q1 vdd 9.49fF
C45 Q0 vdd 5.33fF
C46 DFlipFlop_1/latch_diff_0/m1_657_280# CLK 0.28fF
C47 DFlipFlop_0/Q nCLK 0.11fF
C48 DFlipFlop_0/D sky130_fd_sc_hs__and2_1_0/a_56_136# 0.04fF
C49 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop_1/D 0.03fF
C50 Q1 DFlipFlop_2/nQ 0.31fF
C51 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out nCLK 0.05fF
C52 nCLK vdd 0.34fF
C53 Q1 DFlipFlop_0/latch_diff_1/nD 0.10fF
C54 Q0 DFlipFlop_0/latch_diff_1/nD 0.21fF
C55 sky130_fd_sc_hs__xor2_1_0/a_355_368# vdd 0.03fF
C56 Q1 DFlipFlop_3/nQ 0.10fF
C57 CLK nQ2 0.17fF
C58 sky130_fd_sc_hs__and2_1_1/a_56_136# CLK 0.06fF
C59 DFlipFlop_0/D vdd 0.19fF
C60 sky130_fd_sc_hs__and2_1_0/a_56_136# vdd 0.02fF
C61 nCLK DFlipFlop_2/nQ 0.09fF
C62 Q1 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.09fF
C63 Q0 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.33fF
C64 DFlipFlop_0/latch_diff_1/nD nCLK 0.05fF
C65 Q0 sky130_fd_sc_hs__xor2_1_0/a_194_125# 0.26fF
C66 sky130_fd_sc_hs__or2_1_0/a_63_368# Q1_shift -0.27fF
C67 DFlipFlop_3/nQ nCLK 0.02fF
C68 DFlipFlop_2/D CLK 0.14fF
C69 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vdd 0.03fF
C70 CLK DFlipFlop_3/latch_diff_0/D 0.11fF
C71 CLK_5 vdd 0.15fF
C72 Q1 DFlipFlop_3/latch_diff_0/nD 0.08fF
C73 sky130_fd_sc_hs__xor2_1_0/a_194_125# nCLK 0.11fF
C74 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in CLK 0.03fF
C75 nQ0 CLK 0.19fF
C76 Q1 sky130_fd_sc_hs__and2_1_0/a_143_136# 0.02fF
C77 DFlipFlop_2/nQ vdd 0.02fF
C78 Q0 sky130_fd_sc_hs__and2_1_0/a_143_136# 0.03fF
C79 DFlipFlop_0/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.02fF
C80 DFlipFlop_0/latch_diff_1/m1_657_280# nCLK 0.28fF
C81 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vdd 0.02fF
C82 DFlipFlop_3/latch_diff_0/nD nCLK 0.08fF
C83 nQ0 DFlipFlop_1/latch_diff_1/D 0.91fF
C84 DFlipFlop_0/latch_diff_1/D CLK 0.03fF
C85 DFlipFlop_3/nQ vdd 0.02fF
C86 nQ0 DFlipFlop_1/latch_diff_0/D 0.09fF
C87 Q1 DFlipFlop_2/latch_diff_1/nD 0.21fF
C88 Q1 DFlipFlop_3/latch_diff_1/D 0.79fF
C89 nQ0 DFlipFlop_1/latch_diff_0/nD 0.08fF
C90 CLK DFlipFlop_1/D 0.21fF
C91 sky130_fd_sc_hs__and2_1_1/a_143_136# CLK 0.03fF
C92 sky130_fd_sc_hs__xor2_1_0/a_455_87# DFlipFlop_2/D 0.08fF
C93 DFlipFlop_2/latch_diff_1/D CLK 0.14fF
C94 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vdd 0.02fF
C95 DFlipFlop_1/latch_diff_1/nD CLK 0.09fF
C96 Q1 CLK -0.10fF
C97 sky130_fd_sc_hs__xor2_1_0/a_194_125# vdd 0.03fF
C98 sky130_fd_sc_hs__and2_1_1/a_56_136# nQ2 0.01fF
C99 Q0 CLK 0.08fF
C100 Q1 DFlipFlop_2/latch_diff_1/m1_657_280# 0.03fF
C101 nQ0 DFlipFlop_1/latch_diff_0/m1_657_280# 0.25fF
C102 DFlipFlop_2/latch_diff_1/nD nCLK 0.16fF
C103 DFlipFlop_3/latch_diff_1/D nCLK 0.14fF
C104 Q1 sky130_fd_sc_hs__or2_1_0/a_63_368# 0.10fF
C105 Q1 DFlipFlop_1/latch_diff_1/D -0.10fF
C106 DFlipFlop_1/latch_diff_1/D Q0 0.06fF
C107 Q1 DFlipFlop_1/latch_diff_0/D 0.18fF
C108 Q0 DFlipFlop_1/latch_diff_0/D 0.42fF
C109 Q1 DFlipFlop_2/latch_diff_0/D 0.42fF
C110 DFlipFlop_2/latch_diff_1/m1_657_280# nCLK 0.28fF
C111 Q1 DFlipFlop_3/latch_diff_1/nD 1.24fF
C112 Q1 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in 0.20fF
C113 DFlipFlop_3/latch_diff_1/m1_657_280# Q1 0.28fF
C114 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out CLK -0.31fF
C115 DFlipFlop_1/latch_diff_1/D nCLK 0.08fF
C116 Q1 DFlipFlop_0/latch_diff_0/D 0.15fF
C117 nQ0 nQ2 0.03fF
C118 sky130_fd_sc_hs__and2_1_1/a_56_136# nQ0 0.01fF
C119 Q0 DFlipFlop_0/latch_diff_0/D 0.42fF
C120 DFlipFlop_1/latch_diff_0/D nCLK 0.11fF
C121 DFlipFlop_2/latch_diff_0/D nCLK 0.11fF
C122 DFlipFlop_0/Q CLK 0.08fF
C123 DFlipFlop_3/latch_diff_1/nD nCLK 0.09fF
C124 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in nCLK -0.33fF
C125 CLK vdd 0.41fF
C126 Q1 DFlipFlop_3/latch_diff_0/m1_657_280# 0.28fF
C127 sky130_fd_sc_hs__and2_1_1/a_56_136# DFlipFlop_1/D 0.04fF
C128 sky130_fd_sc_hs__xor2_1_0/a_455_87# nCLK 0.02fF
C129 sky130_fd_sc_hs__and2_1_1/a_143_136# nQ2 0.01fF
C130 Q1 nQ2 0.07fF
C131 Q0 nQ2 0.23fF
C132 Q1 Q1_shift 0.36fF
C133 sky130_fd_sc_hs__or2_1_0/a_63_368# vdd 0.02fF
C134 CLK DFlipFlop_2/nQ 0.13fF
C135 DFlipFlop_3/latch_diff_0/m1_657_280# nCLK 0.27fF
C136 sky130_fd_sc_hs__or2_1_0/a_63_368# CLK_5 0.06fF
C137 CLK DFlipFlop_0/latch_diff_1/nD 0.02fF
C138 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out CLK 0.15fF
C139 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vdd 0.03fF
C140 DFlipFlop_2/D DFlipFlop_1/latch_diff_1/m1_657_280# 0.04fF
C141 Q1 DFlipFlop_2/D 0.10fF
C142 CLK DFlipFlop_3/nQ 0.01fF
C143 nQ2 nCLK 0.10fF
C144 DFlipFlop_2/D Q0 0.25fF
C145 Q1 DFlipFlop_3/latch_diff_0/D 0.09fF
C146 nQ0 DFlipFlop_1/D 0.12fF
C147 sky130_fd_sc_hs__and2_1_1/a_143_136# nQ0 0.04fF
C148 nQ0 DFlipFlop_1/latch_diff_1/m1_657_280# 0.21fF
C149 DFlipFlop_2/latch_diff_0/nD CLK 0.08fF
C150 nQ0 DFlipFlop_1/latch_diff_1/nD 0.88fF
C151 Q1 nQ0 0.06fF
C152 nQ0 Q0 0.33fF
C153 DFlipFlop_2/D nCLK 0.41fF
C154 DFlipFlop_0/Q nQ2 0.09fF
C155 Q1 DFlipFlop_0/latch_diff_1/D 0.06fF
C156 nQ2 vdd 0.04fF
C157 CLK_5 vss -0.18fF
C158 sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.38fF
C159 sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.41fF
C160 sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C161 DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.64fF
C162 Q1_shift vss -0.29fF
C163 DFlipFlop_3/nQ vss 0.52fF
C164 DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C165 DFlipFlop_3/latch_diff_1/D vss -1.73fF
C166 DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C167 DFlipFlop_3/latch_diff_0/D vss 0.96fF
C168 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.94fF
C169 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.64fF
C170 Q1 vss 8.55fF
C171 DFlipFlop_3/latch_diff_0/nD vss 0.94fF
C172 DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.62fF
C173 Q0 vss 0.53fF
C174 nQ0 vss 3.42fF
C175 DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C176 DFlipFlop_1/latch_diff_1/D vss -1.73fF
C177 DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C178 DFlipFlop_1/latch_diff_0/D vss 0.96fF
C179 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C180 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.58fF
C181 DFlipFlop_1/D vss 3.72fF
C182 DFlipFlop_1/latch_diff_0/nD vss 0.94fF
C183 DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.72fF
C184 DFlipFlop_2/nQ vss 0.50fF
C185 DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C186 DFlipFlop_2/latch_diff_1/D vss -1.72fF
C187 DFlipFlop_2/latch_diff_1/nD vss 0.58fF
C188 DFlipFlop_2/latch_diff_0/D vss 0.96fF
C189 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.89fF
C190 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C191 DFlipFlop_2/D vss 5.34fF
C192 DFlipFlop_2/latch_diff_0/nD vss 0.94fF
C193 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.61fF
C194 nCLK vss 0.89fF
C195 DFlipFlop_0/Q vss -0.94fF
C196 nQ2 vss 2.05fF
C197 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C198 CLK vss 0.07fF
C199 DFlipFlop_0/latch_diff_1/D vss -1.73fF
C200 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C201 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C202 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.88fF
C203 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C204 DFlipFlop_0/D vss 4.04fF
C205 vdd vss 144.09fF
C206 DFlipFlop_0/latch_diff_0/nD vss 0.94fF
C207 sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C208 sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.42fF
.ends

.subckt mux2to4 vss out_b_1 vdd select_0 select_0_neg out_a_0 out_a_1 out_b_0 in_a
+ in_b
Xtrans_gate_mux2to8_0 in_a vss out_a_0 select_0_neg select_0 vdd trans_gate_mux2to8
Xtrans_gate_mux2to8_1 in_a vss out_a_1 select_0 select_0_neg vdd trans_gate_mux2to8
Xtrans_gate_mux2to8_2 in_b vss out_b_0 select_0_neg select_0 vdd trans_gate_mux2to8
Xtrans_gate_mux2to8_3 in_b vss out_b_1 select_0 select_0_neg vdd trans_gate_mux2to8
C0 select_0 out_a_1 0.18fF
C1 vdd out_a_1 0.06fF
C2 vdd select_0 0.02fF
C3 select_0_neg in_a 0.22fF
C4 out_b_0 in_a 0.11fF
C5 out_b_0 select_0_neg -0.13fF
C6 in_b select_0_neg 0.10fF
C7 in_b out_b_0 0.08fF
C8 out_a_0 in_a 0.08fF
C9 in_b out_b_1 0.08fF
C10 out_a_0 select_0_neg 0.05fF
C11 out_a_1 in_a 0.08fF
C12 out_a_1 select_0_neg 0.12fF
C13 out_b_0 out_a_1 0.88fF
C14 select_0 in_a 0.31fF
C15 select_0 select_0_neg 0.49fF
C16 select_0 out_b_0 0.03fF
C17 vdd in_a 0.02fF
C18 in_b out_a_1 0.08fF
C19 vdd select_0_neg 0.02fF
C20 vdd out_b_0 0.06fF
C21 in_b select_0 0.24fF
C22 out_b_1 select_0 0.14fF
C23 vdd in_b 0.02fF
C24 vdd out_b_1 0.06fF
C25 vdd out_a_0 0.06fF
C26 out_b_1 vss 0.99fF
C27 in_b vss 2.00fF
C28 out_b_0 vss 0.93fF
C29 out_a_1 vss 0.22fF
C30 vdd vss 9.53fF
C31 in_a vss 2.00fF
C32 out_a_0 vss 0.99fF
C33 select_0_neg vss 2.56fF
C34 select_0 vss 2.23fF
.ends

.subckt sky130_fd_sc_hs__mux2_1 A0 A1 S VGND VNB VPB VPWR X a_304_74# a_443_74# a_524_368#
+ a_27_112#
X0 VPWR S a_27_112# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND a_27_112# a_443_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 X a_304_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VPWR a_27_112# a_524_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_304_74# A1 a_226_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 X a_304_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 a_223_368# S VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_304_74# A0 a_223_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_443_74# A0 a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_524_368# A1 a_304_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_226_74# S VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 VGND S a_27_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
C0 a_524_368# a_27_112# 0.06fF
C1 A1 A0 0.31fF
C2 S A1 0.10fF
C3 VGND A0 0.02fF
C4 VGND S 0.07fF
C5 a_304_74# A0 0.23fF
C6 S a_304_74# 0.18fF
C7 VPWR S 0.05fF
C8 a_27_112# A0 0.07fF
C9 S a_27_112# 0.22fF
C10 VGND A1 0.09fF
C11 X A1 0.02fF
C12 a_304_74# A1 0.69fF
C13 VGND X 0.11fF
C14 VGND a_304_74# 0.58fF
C15 X a_304_74# 0.29fF
C16 VPWR A1 0.01fF
C17 VGND VPWR 0.02fF
C18 a_223_368# a_304_74# 0.05fF
C19 a_443_74# A1 0.07fF
C20 a_304_74# a_226_74# 0.08fF
C21 VPWR X 0.28fF
C22 VPWR VPB 0.06fF
C23 VPWR a_304_74# 0.13fF
C24 a_27_112# A1 0.18fF
C25 VGND a_27_112# 0.18fF
C26 a_443_74# a_304_74# 0.12fF
C27 X a_27_112# 0.08fF
C28 a_27_112# VPB 0.01fF
C29 a_304_74# a_27_112# 0.58fF
C30 a_223_368# a_27_112# 0.09fF
C31 S A0 0.04fF
C32 VPWR a_27_112# 0.99fF
C33 VGND VNB 0.88fF
C34 X VNB 0.25fF
C35 VPWR VNB 0.89fF
C36 A1 VNB 0.37fF
C37 A0 VNB 0.23fF
C38 S VNB 0.34fF
C39 VPB VNB 0.87fF
C40 a_304_74# VNB 0.36fF
C41 a_27_112# VNB 0.65fF
.ends

.subckt prescaler_23 nCLK vss DFlipFlop_0/latch_diff_1/nD nCLK_23 DFlipFlop_2/latch_diff_0/nD
+ vdd DFlipFlop_2/latch_diff_1/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out CLK_23 DFlipFlop_2/latch_diff_0/m1_657_280#
+ DFlipFlop_0/latch_diff_0/D CLK DFlipFlop_2/latch_diff_1/nD DFlipFlop_2/latch_diff_1/m1_657_280#
+ DFlipFlop_0/latch_diff_1/D DFlipFlop_0/latch_diff_0/nD MC DFlipFlop_2/latch_diff_0/D
+ Q2
Xsky130_fd_sc_hs__mux2_1_0 sky130_fd_sc_hs__or2_1_1/X nCLK_23 MC vss vss vdd vdd CLK_23
+ sky130_fd_sc_hs__mux2_1_0/a_304_74# sky130_fd_sc_hs__mux2_1_0/a_443_74# sky130_fd_sc_hs__mux2_1_0/a_524_368#
+ sky130_fd_sc_hs__mux2_1_0/a_27_112# sky130_fd_sc_hs__mux2_1
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vdd vss DFlipFlop_0/latch_diff_1/D
+ DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_0/nQ nCLK DFlipFlop_0/latch_diff_0/nD
+ Q1 DFlipFlop_0/latch_diff_1/nD nCLK_23 DFlipFlop_0/latch_diff_1/m1_657_280# DFlipFlop_0/latch_diff_0/D
+ CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop
XDFlipFlop_1 DFlipFlop_1/latch_diff_0/m1_657_280# vdd vss DFlipFlop_1/latch_diff_1/D
+ DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in nCLK_23 nCLK DFlipFlop_1/latch_diff_0/nD
+ Q2 DFlipFlop_1/latch_diff_1/nD DFlipFlop_1/D DFlipFlop_1/latch_diff_1/m1_657_280#
+ DFlipFlop_1/latch_diff_0/D CLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop
XDFlipFlop_2 DFlipFlop_2/latch_diff_0/m1_657_280# vdd vss DFlipFlop_2/latch_diff_1/D
+ DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_2/nQ CLK DFlipFlop_2/latch_diff_0/nD
+ Q2_d DFlipFlop_2/latch_diff_1/nD Q2 DFlipFlop_2/latch_diff_1/m1_657_280# DFlipFlop_2/latch_diff_0/D
+ nCLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop
Xsky130_fd_sc_hs__and2_1_0 nCLK_23 sky130_fd_sc_hs__or2_1_0/X vss vss vdd vdd DFlipFlop_1/D
+ sky130_fd_sc_hs__and2_1_0/a_143_136# sky130_fd_sc_hs__and2_1_0/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__or2_1_0 Q1 MC vss vss vdd vdd sky130_fd_sc_hs__or2_1_0/X sky130_fd_sc_hs__or2_1_0/a_152_368#
+ sky130_fd_sc_hs__or2_1_0/a_63_368# sky130_fd_sc_hs__or2_1
Xsky130_fd_sc_hs__or2_1_1 Q2 Q2_d vss vss vdd vdd sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__or2_1_1/a_152_368#
+ sky130_fd_sc_hs__or2_1_1/a_63_368# sky130_fd_sc_hs__or2_1
C0 nCLK vdd -0.55fF
C1 DFlipFlop_2/nQ CLK 0.02fF
C2 CLK sky130_fd_sc_hs__or2_1_0/X 0.01fF
C3 Q1 MC 0.29fF
C4 sky130_fd_sc_hs__mux2_1_0/a_27_112# MC 0.24fF
C5 CLK DFlipFlop_1/D 0.40fF
C6 DFlipFlop_2/latch_diff_1/D Q2 0.13fF
C7 sky130_fd_sc_hs__and2_1_0/a_56_136# CLK 0.08fF
C8 DFlipFlop_1/latch_diff_0/nD CLK 0.09fF
C9 DFlipFlop_2/latch_diff_1/D CLK 0.09fF
C10 Q2 sky130_fd_sc_hs__or2_1_1/X 0.24fF
C11 DFlipFlop_2/nQ nCLK 0.02fF
C12 nCLK sky130_fd_sc_hs__or2_1_0/X 0.06fF
C13 nCLK DFlipFlop_1/D 0.16fF
C14 DFlipFlop_0/latch_diff_0/m1_657_280# CLK 0.29fF
C15 sky130_fd_sc_hs__or2_1_1/a_63_368# Q2 0.09fF
C16 nCLK DFlipFlop_2/latch_diff_1/D 0.16fF
C17 DFlipFlop_2/latch_diff_1/m1_657_280# CLK 0.33fF
C18 sky130_fd_sc_hs__mux2_1_0/a_443_74# nCLK_23 0.09fF
C19 vdd nCLK_23 3.27fF
C20 nCLK sky130_fd_sc_hs__or2_1_0/a_152_368# 0.01fF
C21 CLK DFlipFlop_1/latch_diff_0/m1_657_280# 0.31fF
C22 nCLK DFlipFlop_1/latch_diff_1/m1_657_280# 0.31fF
C23 sky130_fd_sc_hs__or2_1_0/a_63_368# Q1 0.09fF
C24 nCLK_23 sky130_fd_sc_hs__or2_1_0/X 0.07fF
C25 CLK Q2 0.29fF
C26 DFlipFlop_1/latch_diff_1/D CLK 0.18fF
C27 nCLK_23 DFlipFlop_1/D 0.02fF
C28 sky130_fd_sc_hs__and2_1_0/a_56_136# nCLK_23 0.14fF
C29 vdd Q1 0.07fF
C30 nCLK_23 DFlipFlop_0/latch_diff_0/nD 0.12fF
C31 sky130_fd_sc_hs__mux2_1_0/a_524_368# nCLK_23 0.04fF
C32 nCLK Q2 0.29fF
C33 nCLK DFlipFlop_1/latch_diff_1/D 0.09fF
C34 CLK DFlipFlop_0/latch_diff_1/nD 0.02fF
C35 nCLK_23 sky130_fd_sc_hs__or2_1_1/X 0.26fF
C36 vdd DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out 0.03fF
C37 Q1 sky130_fd_sc_hs__or2_1_0/X 0.06fF
C38 vdd MC 0.88fF
C39 DFlipFlop_1/latch_diff_1/nD CLK 0.11fF
C40 nCLK DFlipFlop_0/latch_diff_1/nD 0.05fF
C41 nCLK DFlipFlop_0/latch_diff_1/m1_657_280# 0.28fF
C42 DFlipFlop_2/latch_diff_0/D Q2 0.30fF
C43 sky130_fd_sc_hs__or2_1_0/X MC 0.09fF
C44 sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__mux2_1_0/a_304_74# 0.08fF
C45 DFlipFlop_2/latch_diff_0/D CLK 0.13fF
C46 nCLK DFlipFlop_1/latch_diff_1/nD 0.18fF
C47 Q1 sky130_fd_sc_hs__or2_1_0/a_152_368# 0.01fF
C48 nCLK_23 Q2 0.03fF
C49 nCLK_23 CLK 0.22fF
C50 sky130_fd_sc_hs__or2_1_1/X MC 0.02fF
C51 vdd DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in 0.03fF
C52 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out CLK 0.16fF
C53 nCLK_23 DFlipFlop_0/latch_diff_1/nD 0.02fF
C54 DFlipFlop_0/latch_diff_1/D CLK 0.04fF
C55 nCLK nCLK_23 0.11fF
C56 Q1 CLK -0.07fF
C57 DFlipFlop_0/nQ CLK 0.15fF
C58 CLK_23 sky130_fd_sc_hs__mux2_1_0/a_304_74# 0.05fF
C59 Q1 DFlipFlop_0/latch_diff_1/nD 0.03fF
C60 vdd Q2_d 0.02fF
C61 Q2 MC 0.18fF
C62 DFlipFlop_0/latch_diff_1/m1_657_280# Q1 0.06fF
C63 nCLK Q1 -0.02fF
C64 nCLK DFlipFlop_0/nQ 0.11fF
C65 DFlipFlop_2/latch_diff_1/nD Q2 0.17fF
C66 nCLK_23 sky130_fd_sc_hs__and2_1_0/a_143_136# 0.02fF
C67 vdd sky130_fd_sc_hs__or2_1_0/X 0.03fF
C68 CLK MC 0.08fF
C69 vdd DFlipFlop_1/D 0.07fF
C70 DFlipFlop_2/latch_diff_1/nD CLK 0.19fF
C71 nCLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out 0.06fF
C72 nCLK DFlipFlop_2/latch_diff_0/m1_657_280# 0.31fF
C73 nCLK MC 0.01fF
C74 sky130_fd_sc_hs__mux2_1_0/a_443_74# sky130_fd_sc_hs__or2_1_1/X 0.03fF
C75 DFlipFlop_0/latch_diff_1/D nCLK_23 0.05fF
C76 DFlipFlop_2/latch_diff_1/D Q2_d 0.03fF
C77 sky130_fd_sc_hs__or2_1_0/X DFlipFlop_1/D 0.35fF
C78 vdd sky130_fd_sc_hs__or2_1_1/X 0.03fF
C79 DFlipFlop_2/latch_diff_1/nD nCLK 0.12fF
C80 nCLK_23 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.49fF
C81 sky130_fd_sc_hs__and2_1_0/a_56_136# sky130_fd_sc_hs__or2_1_0/X 0.07fF
C82 Q2_d sky130_fd_sc_hs__or2_1_1/X 0.03fF
C83 nCLK DFlipFlop_2/latch_diff_0/nD 0.09fF
C84 nCLK_23 Q1 0.02fF
C85 Q2 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in 0.38fF
C86 nCLK_23 DFlipFlop_0/nQ 0.05fF
C87 nCLK_23 sky130_fd_sc_hs__mux2_1_0/a_304_74# 0.04fF
C88 sky130_fd_sc_hs__mux2_1_0/a_27_112# nCLK_23 0.07fF
C89 DFlipFlop_2/latch_diff_1/m1_657_280# Q2_d 0.03fF
C90 nCLK DFlipFlop_1/latch_diff_0/D 0.02fF
C91 CLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in -0.10fF
C92 nCLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in -0.02fF
C93 nCLK_23 MC 4.46fF
C94 vdd Q2 1.63fF
C95 DFlipFlop_0/nQ Q1 -0.02fF
C96 Q2_d Q2 0.66fF
C97 vdd CLK 0.34fF
C98 nCLK sky130_fd_sc_hs__or2_1_0/a_63_368# 0.05fF
C99 CLK_23 vdd 0.16fF
C100 DFlipFlop_2/nQ Q2 0.13fF
C101 sky130_fd_sc_hs__or2_1_1/a_63_368# vss 0.37fF
C102 sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C103 sky130_fd_sc_hs__or2_1_0/X vss 0.92fF
C104 sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.39fF
C105 DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C106 Q2_d vss -0.22fF
C107 DFlipFlop_2/nQ vss 0.48fF
C108 DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C109 DFlipFlop_2/latch_diff_1/D vss -1.73fF
C110 DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C111 DFlipFlop_2/latch_diff_0/D vss 0.96fF
C112 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.94fF
C113 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.63fF
C114 Q2 vss 1.35fF
C115 DFlipFlop_2/latch_diff_0/nD vss 0.94fF
C116 DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.72fF
C117 DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C118 DFlipFlop_1/latch_diff_1/D vss -1.72fF
C119 DFlipFlop_1/latch_diff_1/nD vss 0.58fF
C120 DFlipFlop_1/latch_diff_0/D vss 0.96fF
C121 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C122 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C123 DFlipFlop_1/D vss 2.98fF
C124 DFlipFlop_1/latch_diff_0/nD vss 0.94fF
C125 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C126 nCLK vss -1.56fF
C127 Q1 vss 0.50fF
C128 DFlipFlop_0/nQ vss 0.48fF
C129 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C130 CLK vss -0.69fF
C131 DFlipFlop_0/latch_diff_1/D vss -1.73fF
C132 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C133 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C134 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C135 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C136 nCLK_23 vss -0.65fF
C137 vdd vss 113.67fF
C138 DFlipFlop_0/latch_diff_0/nD vss 0.94fF
C139 CLK_23 vss -0.57fF
C140 sky130_fd_sc_hs__or2_1_1/X vss -0.35fF
C141 MC vss 2.09fF
C142 sky130_fd_sc_hs__mux2_1_0/a_304_74# vss 0.41fF
C143 sky130_fd_sc_hs__mux2_1_0/a_27_112# vss 0.69fF
.ends

.subckt freq_div clk_0 vss n_clk_0 vdd prescaler_23_0/Q2 s_0 s_1_n s_1 prescaler_23_0/nCLK_23
+ prescaler_23_0/MC clk_d prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# s_0_n
+ clk_pre div_by_5_0/DFlipFlop_2/latch_diff_0/nD prescaler_23_0/DFlipFlop_2/latch_diff_1/D
+ prescaler_23_0/DFlipFlop_2/latch_diff_1/nD clk_1 div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280#
+ clk_out_mux21 n_clk_1 out div_by_5_0/Q1 div_by_5_0/DFlipFlop_2/latch_diff_0/D prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280#
+ div_by_5_0/DFlipFlop_2/latch_diff_1/nD clk_2 in_a in_b clk_5 prescaler_23_0/DFlipFlop_2/latch_diff_0/D
+ prescaler_23_0/DFlipFlop_2/latch_diff_0/nD div_by_5_0/DFlipFlop_2/latch_diff_1/D
Xdiv_by_2_0 vdd vss div_by_2_0/nout_div clk_2 div_by_2_0/nCLK_2 div_by_2_0/o1 div_by_2_0/o2
+ clk_out_mux21 div_by_2_0/out_div div_by_2
Xmux2to1_0 vss s_0_n clk_pre clk_5 s_0 vdd clk_out_mux21 mux2to1
Xinverter_min_x4_0 inverter_min_x4_0/in vss clk_d vdd inverter_min_x4
Xmux2to1_1 vss s_1_n clk_d clk_2 s_1 vdd out mux2to1
Xinverter_min_x2_0 clk_out_mux21 inverter_min_x4_0/in vss vdd inverter_min_x2
Xinverter_min_x2_1 s_1 s_1_n vss vdd inverter_min_x2
Xinverter_min_x2_2 s_0 s_0_n vss vdd inverter_min_x2
Xdiv_by_5_0 n_clk_1 div_by_5_0/DFlipFlop_0/latch_diff_1/nD div_by_5_0/DFlipFlop_2/latch_diff_0/nD
+ vss div_by_5_0/Q1 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in clk_1
+ div_by_5_0/DFlipFlop_0/Q vdd div_by_5_0/DFlipFlop_2/latch_diff_1/D div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# div_by_5_0/DFlipFlop_3/latch_diff_0/D
+ div_by_5_0/DFlipFlop_3/latch_diff_1/nD div_by_5_0/DFlipFlop_1/latch_diff_1/nD div_by_5_0/DFlipFlop_1/latch_diff_0/nD
+ div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# clk_5 div_by_5_0/Q1_shift div_by_5_0/nQ2
+ div_by_5_0/DFlipFlop_0/latch_diff_0/D div_by_5_0/DFlipFlop_2/D div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_1/latch_diff_1/D div_by_5_0/DFlipFlop_1/D div_by_5_0/nQ0 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ div_by_5_0/DFlipFlop_2/latch_diff_1/nD div_by_5_0/Q0 div_by_5_0/DFlipFlop_0/D div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_0/latch_diff_1/D div_by_5_0/DFlipFlop_0/latch_diff_0/nD div_by_5_0/DFlipFlop_2/nQ
+ div_by_5_0/DFlipFlop_2/latch_diff_0/D div_by_5_0/DFlipFlop_3/latch_diff_1/D div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_152_368#
+ div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# div_by_5_0/DFlipFlop_3/nQ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136#
+ div_by_5
Xmux2to4_0 vss n_clk_1 vdd s_0 s_0_n clk_0 clk_1 n_clk_0 in_a in_b mux2to4
Xprescaler_23_0 n_clk_0 vss prescaler_23_0/DFlipFlop_0/latch_diff_1/nD prescaler_23_0/nCLK_23
+ prescaler_23_0/DFlipFlop_2/latch_diff_0/nD vdd prescaler_23_0/DFlipFlop_2/latch_diff_1/D
+ prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ clk_pre prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# prescaler_23_0/DFlipFlop_0/latch_diff_0/D
+ clk_0 prescaler_23_0/DFlipFlop_2/latch_diff_1/nD prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280#
+ prescaler_23_0/DFlipFlop_0/latch_diff_1/D prescaler_23_0/DFlipFlop_0/latch_diff_0/nD
+ prescaler_23_0/MC prescaler_23_0/DFlipFlop_2/latch_diff_0/D prescaler_23_0/Q2 prescaler_23
C0 s_0 div_by_5_0/DFlipFlop_3/latch_diff_1/nD 0.05fF
C1 div_by_5_0/DFlipFlop_2/latch_diff_1/D s_0_n 0.04fF
C2 clk_0 vdd 0.63fF
C3 s_0_n div_by_5_0/DFlipFlop_2/latch_diff_1/nD 0.24fF
C4 s_0 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out -0.13fF
C5 clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_1/nD 0.09fF
C6 vdd s_0_n 2.53fF
C7 div_by_5_0/DFlipFlop_0/D s_0_n 0.05fF
C8 div_by_5_0/Q0 s_0 0.02fF
C9 s_0 div_by_5_0/DFlipFlop_2/D 0.03fF
C10 s_0 clk_out_mux21 0.68fF
C11 n_clk_0 prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.14fF
C12 out s_1 0.39fF
C13 s_0 div_by_5_0/DFlipFlop_1/latch_diff_1/D 0.05fF
C14 s_0 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out -0.19fF
C15 s_1_n clk_2 0.59fF
C16 s_0 div_by_5_0/DFlipFlop_2/latch_diff_0/nD 0.12fF
C17 s_0 clk_pre 0.21fF
C18 vdd n_clk_1 0.13fF
C19 div_by_5_0/DFlipFlop_0/D n_clk_1 0.21fF
C20 in_a s_0 0.30fF
C21 clk_1 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.08fF
C22 s_0_n div_by_5_0/DFlipFlop_3/latch_diff_1/D 0.24fF
C23 n_clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_1/D 0.09fF
C24 clk_5 s_0_n 0.56fF
C25 n_clk_0 clk_1 -0.03fF
C26 s_0 div_by_5_0/DFlipFlop_1/latch_diff_1/nD 0.02fF
C27 clk_pre clk_out_mux21 1.19fF
C28 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in n_clk_1 0.14fF
C29 s_0 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in -0.36fF
C30 clk_d inverter_min_x4_0/in 0.11fF
C31 s_0 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out 0.30fF
C32 div_by_5_0/Q1_shift s_0_n 0.04fF
C33 n_clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_0/D 0.13fF
C34 s_0 clk_1 1.36fF
C35 s_0 div_by_5_0/DFlipFlop_1/D 0.03fF
C36 s_0 div_by_5_0/DFlipFlop_0/latch_diff_1/D 0.05fF
C37 clk_1 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out 0.05fF
C38 prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out clk_0 0.16fF
C39 s_0 div_by_5_0/nQ0 0.05fF
C40 s_0 div_by_5_0/DFlipFlop_3/latch_diff_0/D 0.10fF
C41 s_0_n div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.24fF
C42 n_clk_0 s_0_n 0.31fF
C43 s_0 div_by_5_0/nQ2 0.05fF
C44 clk_5 vdd 0.04fF
C45 div_by_5_0/DFlipFlop_3/nQ s_0 0.02fF
C46 div_by_5_0/DFlipFlop_2/nQ s_0_n 0.04fF
C47 s_0 div_by_5_0/DFlipFlop_1/latch_diff_0/nD 0.12fF
C48 s_0_n div_by_5_0/DFlipFlop_0/Q 0.24fF
C49 out clk_2 0.05fF
C50 n_clk_1 div_by_5_0/DFlipFlop_0/latch_diff_0/D 0.11fF
C51 s_0 s_0_n 7.76fF
C52 s_0_n div_by_5_0/Q1 0.21fF
C53 div_by_5_0/DFlipFlop_3/latch_diff_1/nD s_0_n 0.04fF
C54 n_clk_0 prescaler_23_0/nCLK_23 0.16fF
C55 s_0 div_by_5_0/DFlipFlop_0/latch_diff_0/nD 0.12fF
C56 n_clk_1 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.11fF
C57 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out s_0_n -0.01fF
C58 in_a clk_1 0.05fF
C59 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# n_clk_1 0.06fF
C60 div_by_5_0/Q0 s_0_n 0.24fF
C61 s_0_n div_by_5_0/DFlipFlop_2/D 0.05fF
C62 vdd clk_2 0.02fF
C63 n_clk_0 vdd 0.25fF
C64 clk_out_mux21 s_0_n 0.45fF
C65 n_clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_1/nD 0.13fF
C66 div_by_5_0/Q1_shift div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_152_368# -0.02fF
C67 s_0 div_by_5_0/DFlipFlop_2/latch_diff_1/D 0.05fF
C68 n_clk_1 div_by_5_0/Q1 0.15fF
C69 div_by_5_0/DFlipFlop_1/latch_diff_1/D s_0_n 0.04fF
C70 s_0 div_by_5_0/DFlipFlop_2/latch_diff_1/nD 0.02fF
C71 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out s_0_n -0.29fF
C72 div_by_5_0/DFlipFlop_2/latch_diff_0/nD s_0_n 0.20fF
C73 s_0 vdd 3.67fF
C74 vdd div_by_5_0/Q1 -0.02fF
C75 div_by_5_0/DFlipFlop_0/D s_0 0.03fF
C76 div_by_5_0/DFlipFlop_0/D div_by_5_0/Q1 -0.02fF
C77 clk_5 div_by_5_0/Q1_shift 0.04fF
C78 div_by_5_0/Q0 n_clk_1 0.01fF
C79 in_b s_0_n 0.48fF
C80 clk_1 div_by_5_0/DFlipFlop_0/latch_diff_1/D 0.11fF
C81 div_by_5_0/Q0 vdd 0.05fF
C82 clk_pre prescaler_23_0/nCLK_23 0.03fF
C83 div_by_5_0/DFlipFlop_1/latch_diff_1/nD s_0_n 0.24fF
C84 vdd clk_out_mux21 0.14fF
C85 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/Q1 -0.06fF
C86 clk_d s_1 0.22fF
C87 clk_d vdd 0.23fF
C88 prescaler_23_0/DFlipFlop_0/latch_diff_1/D clk_0 0.13fF
C89 out s_1_n 0.33fF
C90 s_0_n div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in -0.37fF
C91 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out s_0_n 0.31fF
C92 clk_1 s_0_n 4.82fF
C93 in_b n_clk_1 0.05fF
C94 clk_pre vdd 0.17fF
C95 div_by_5_0/DFlipFlop_1/D s_0_n 0.19fF
C96 s_0 div_by_5_0/DFlipFlop_3/latch_diff_1/D 0.02fF
C97 clk_1 div_by_5_0/DFlipFlop_0/latch_diff_0/nD 0.08fF
C98 div_by_5_0/DFlipFlop_0/latch_diff_1/D s_0_n 0.04fF
C99 vdd inverter_min_x4_0/in 0.09fF
C100 div_by_5_0/nQ0 s_0_n 0.05fF
C101 div_by_5_0/DFlipFlop_3/latch_diff_0/D s_0_n 0.17fF
C102 clk_0 prescaler_23_0/DFlipFlop_0/latch_diff_0/nD 0.09fF
C103 s_1_n s_1 0.39fF
C104 s_0_n div_by_5_0/nQ2 0.05fF
C105 div_by_5_0/Q1_shift s_0 0.05fF
C106 div_by_5_0/DFlipFlop_3/nQ s_0_n 0.24fF
C107 s_0_n div_by_5_0/DFlipFlop_1/latch_diff_0/nD 0.20fF
C108 clk_5 clk_out_mux21 0.05fF
C109 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# n_clk_1 0.03fF
C110 clk_1 vdd 0.16fF
C111 n_clk_1 div_by_5_0/DFlipFlop_0/latch_diff_1/D 0.08fF
C112 s_0 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.02fF
C113 div_by_5_0/DFlipFlop_0/D clk_1 0.14fF
C114 s_0_n div_by_5_0/DFlipFlop_0/latch_diff_0/nD 0.20fF
C115 clk_0 prescaler_23_0/nCLK_23 0.16fF
C116 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# s_0_n 0.05fF
C117 s_0 div_by_5_0/DFlipFlop_2/nQ 0.05fF
C118 s_0 div_by_5_0/DFlipFlop_0/Q 0.02fF
C119 s_0 div_by_5_0/Q1 0.04fF
C120 prescaler_23_0/sky130_fd_sc_hs__or2_1_1/a_63_368# vss 0.37fF
C121 prescaler_23_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C122 prescaler_23_0/sky130_fd_sc_hs__or2_1_0/X vss 0.49fF
C123 prescaler_23_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C124 prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C125 prescaler_23_0/Q2_d vss -0.69fF
C126 prescaler_23_0/DFlipFlop_2/nQ vss 0.48fF
C127 prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C128 prescaler_23_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C129 prescaler_23_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C130 prescaler_23_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C131 prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C132 prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C133 prescaler_23_0/Q2 vss 0.55fF
C134 prescaler_23_0/DFlipFlop_2/latch_diff_0/nD vss 0.94fF
C135 prescaler_23_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C136 prescaler_23_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C137 prescaler_23_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C138 prescaler_23_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C139 prescaler_23_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C140 prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C141 prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C142 prescaler_23_0/DFlipFlop_1/D vss 1.90fF
C143 prescaler_23_0/DFlipFlop_1/latch_diff_0/nD vss 0.94fF
C144 prescaler_23_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C145 n_clk_0 vss -5.35fF
C146 prescaler_23_0/Q1 vss 0.07fF
C147 prescaler_23_0/DFlipFlop_0/nQ vss 0.48fF
C148 prescaler_23_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C149 clk_0 vss 0.66fF
C150 prescaler_23_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C151 prescaler_23_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C152 prescaler_23_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C153 prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C154 prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C155 prescaler_23_0/nCLK_23 vss -1.02fF
C156 prescaler_23_0/DFlipFlop_0/latch_diff_0/nD vss 0.94fF
C157 prescaler_23_0/sky130_fd_sc_hs__or2_1_1/X vss -1.01fF
C158 prescaler_23_0/MC vss 1.07fF
C159 prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_304_74# vss 0.36fF
C160 prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_27_112# vss 0.65fF
C161 in_b vss 2.02fF
C162 in_a vss 2.01fF
C163 s_0_n vss -2.51fF
C164 s_0 vss 5.84fF
C165 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C166 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.38fF
C167 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C168 div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.57fF
C169 div_by_5_0/Q1_shift vss -0.36fF
C170 div_by_5_0/DFlipFlop_3/nQ vss 0.48fF
C171 div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C172 div_by_5_0/DFlipFlop_3/latch_diff_1/D vss -1.73fF
C173 div_by_5_0/DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C174 div_by_5_0/DFlipFlop_3/latch_diff_0/D vss 0.96fF
C175 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C176 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C177 div_by_5_0/Q1 vss 4.35fF
C178 div_by_5_0/DFlipFlop_3/latch_diff_0/nD vss 0.94fF
C179 div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C180 div_by_5_0/Q0 vss 0.29fF
C181 div_by_5_0/nQ0 vss 0.99fF
C182 div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C183 div_by_5_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C184 div_by_5_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C185 div_by_5_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C186 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C187 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C188 div_by_5_0/DFlipFlop_1/D vss 3.64fF
C189 div_by_5_0/DFlipFlop_1/latch_diff_0/nD vss 0.94fF
C190 div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C191 div_by_5_0/DFlipFlop_2/nQ vss 0.48fF
C192 div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C193 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C194 div_by_5_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C195 div_by_5_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C196 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C197 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C198 div_by_5_0/DFlipFlop_2/D vss 3.13fF
C199 div_by_5_0/DFlipFlop_2/latch_diff_0/nD vss 0.94fF
C200 div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C201 n_clk_1 vss -0.55fF
C202 div_by_5_0/DFlipFlop_0/Q vss -0.94fF
C203 div_by_5_0/nQ2 vss 1.38fF
C204 div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C205 clk_1 vss -1.34fF
C206 div_by_5_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C207 div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C208 div_by_5_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C209 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C210 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C211 div_by_5_0/DFlipFlop_0/D vss 3.96fF
C212 vdd vss 344.01fF
C213 div_by_5_0/DFlipFlop_0/latch_diff_0/nD vss 0.94fF
C214 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C215 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.40fF
C216 out vss 0.93fF
C217 clk_d vss 0.78fF
C218 s_1_n vss 1.22fF
C219 s_1 vss 2.97fF
C220 inverter_min_x4_0/in vss 2.77fF
C221 clk_out_mux21 vss 5.29fF
C222 clk_pre vss 1.30fF
C223 clk_2 vss 3.46fF
C224 div_by_2_0/o1 vss 2.20fF
C225 div_by_2_0/nCLK_2 vss 1.04fF
C226 div_by_2_0/o2 vss 2.08fF
C227 div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C228 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C229 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C230 div_by_2_0/DFlipFlop_0/nCLK vss 0.82fF
C231 div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C232 div_by_2_0/out_div vss -0.80fF
C233 div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C234 div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C235 div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C236 div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C237 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C238 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C239 div_by_2_0/nout_div vss 2.62fF
C240 div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 0.94fF
.ends

.subckt sky130_fd_pr__pfet_01v8_58ZKDE VSUBS a_n257_n777# a_n129_n600# a_n221_n600#
+ w_n257_n702#
X0 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X1 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X2 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X3 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
C0 a_n257_n777# a_n221_n600# 0.25fF
C1 a_n221_n600# a_n129_n600# 7.87fF
C2 a_n257_n777# a_n129_n600# 0.29fF
C3 a_n129_n600# VSUBS 0.10fF
C4 a_n221_n600# VSUBS 0.25fF
C5 a_n257_n777# VSUBS 1.05fF
C6 w_n257_n702# VSUBS 2.16fF
.ends

.subckt sky130_fd_pr__nfet_01v8_T69Y3A a_n129_n300# a_n221_n300# w_n257_n327# a_n257_n404#
X0 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
C0 a_n221_n300# a_n129_n300# 4.05fF
C1 a_n221_n300# a_n257_n404# 0.21fF
C2 a_n129_n300# a_n257_n404# 0.30fF
C3 a_n129_n300# w_n257_n327# 0.11fF
C4 a_n221_n300# w_n257_n327# 0.25fF
C5 a_n257_n404# w_n257_n327# 1.11fF
.ends

.subckt buffer_salida a_678_n100# out vdd in vss
Xsky130_fd_pr__pfet_01v8_58ZKDE_1 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_2 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_3 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_0 a_678_n100# vss vss in sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_1 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_4 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_5 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_2 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_3 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_6 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_4 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_7 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_70 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_8 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_5 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_71 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_60 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_6 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_9 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_72 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_61 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_50 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_7 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_62 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_51 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_40 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_8 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_63 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_52 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_41 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_30 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_9 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_20 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_64 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_53 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_42 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_31 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_10 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_21 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_65 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_54 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_43 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_32 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_11 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_22 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_66 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_55 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_44 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_33 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_12 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_23 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_67 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_56 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_45 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_34 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_13 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_24 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_68 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_57 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_46 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_35 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_14 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_69 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_58 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_47 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_36 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_25 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_15 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_59 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_48 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_37 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_26 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_16 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_49 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_38 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_27 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_70 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_17 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_39 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_28 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_71 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_60 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_18 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_29 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_72 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_61 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_50 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_19 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_62 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_51 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_40 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_63 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_52 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_41 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_30 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_20 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_64 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_53 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_42 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_31 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_10 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_21 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_65 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_54 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_43 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_32 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_11 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_22 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_66 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_55 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_44 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_33 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_12 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_23 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_67 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_56 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_45 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_34 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_13 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_24 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_68 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_57 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_46 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_35 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_14 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_69 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_58 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_47 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_36 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_25 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_15 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_59 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_48 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_37 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_26 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_16 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_49 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_38 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_27 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_17 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_39 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_28 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_18 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_29 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_19 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_0 vss in a_678_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
C0 vdd in 0.02fF
C1 in a_678_n100# 0.81fF
C2 vdd a_3996_n100# 3.68fF
C3 a_3996_n100# a_678_n100# 6.52fF
C4 vdd a_678_n100# 0.08fF
C5 a_3996_n100# out 55.19fF
C6 vdd out 47.17fF
C7 vdd vss 20.93fF
C8 out vss 35.17fF
C9 a_3996_n100# vss 49.53fF
C10 a_678_n100# vss 13.08fF
C11 in vss 0.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_CBAU6Y a_n73_n150# a_n33_n238# w_n211_n360# a_15_n150#
X0 a_15_n150# a_n33_n238# a_n73_n150# w_n211_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n33_n238# a_15_n150# 0.02fF
C1 a_n73_n150# a_15_n150# 0.51fF
C2 a_n73_n150# a_n33_n238# 0.02fF
C3 a_15_n150# w_n211_n360# 0.23fF
C4 a_n73_n150# w_n211_n360# 0.23fF
C5 a_n33_n238# w_n211_n360# 0.17fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4757AC VSUBS a_n73_n150# a_n33_181# w_n211_n369# a_15_n150#
X0 a_15_n150# a_n33_181# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_15_n150# a_n33_181# 0.01fF
C1 w_n211_n369# a_n73_n150# 0.20fF
C2 a_n33_181# a_n73_n150# 0.01fF
C3 a_n33_181# w_n211_n369# 0.05fF
C4 a_15_n150# a_n73_n150# 0.51fF
C5 a_15_n150# w_n211_n369# 0.20fF
C6 a_15_n150# VSUBS 0.03fF
C7 a_n73_n150# VSUBS 0.03fF
C8 a_n33_181# VSUBS 0.13fF
C9 w_n211_n369# VSUBS 1.98fF
.ends

.subckt sky130_fd_pr__nfet_01v8_7H8F5S a_n465_172# a_n417_n150# a_351_n150# a_255_n150#
+ w_n647_n360# a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150#
X0 a_159_n150# a_n465_172# a_63_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n225_n150# a_n465_172# a_n321_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_447_n150# a_n465_172# a_351_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_63_n150# a_n465_172# a_n33_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n465_172# a_n225_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n465_172# a_n509_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n33_n150# a_n465_172# a_n129_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_351_n150# a_n465_172# a_255_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_255_n150# a_n465_172# a_159_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n321_n150# a_n465_172# a_n417_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_159_n150# a_447_n150# 0.10fF
C1 a_n129_n150# a_255_n150# 0.07fF
C2 a_n129_n150# a_n465_172# 0.10fF
C3 a_n225_n150# a_n321_n150# 0.43fF
C4 a_n321_n150# a_n509_n150# 0.16fF
C5 a_159_n150# a_n33_n150# 0.16fF
C6 a_n225_n150# a_n129_n150# 0.43fF
C7 a_n129_n150# a_n509_n150# 0.07fF
C8 a_351_n150# a_447_n150# 0.43fF
C9 a_447_n150# a_63_n150# 0.07fF
C10 a_351_n150# a_n33_n150# 0.07fF
C11 a_63_n150# a_n33_n150# 0.43fF
C12 a_n465_172# a_n417_n150# 0.10fF
C13 a_n225_n150# a_n417_n150# 0.16fF
C14 a_n509_n150# a_n417_n150# 0.43fF
C15 a_n321_n150# a_n33_n150# 0.10fF
C16 a_n129_n150# a_n33_n150# 0.43fF
C17 a_159_n150# a_351_n150# 0.16fF
C18 a_159_n150# a_63_n150# 0.43fF
C19 a_n33_n150# a_n417_n150# 0.07fF
C20 a_351_n150# a_63_n150# 0.10fF
C21 a_n465_172# a_255_n150# 0.10fF
C22 a_159_n150# a_n129_n150# 0.10fF
C23 a_n225_n150# a_n465_172# 0.10fF
C24 a_n509_n150# a_n465_172# 0.01fF
C25 a_n225_n150# a_n509_n150# 0.10fF
C26 a_n321_n150# a_63_n150# 0.07fF
C27 a_n129_n150# a_63_n150# 0.16fF
C28 a_n129_n150# a_n321_n150# 0.16fF
C29 a_447_n150# a_255_n150# 0.16fF
C30 a_447_n150# a_n465_172# 0.01fF
C31 a_n33_n150# a_255_n150# 0.10fF
C32 a_n33_n150# a_n465_172# 0.10fF
C33 a_n225_n150# a_n33_n150# 0.16fF
C34 a_n321_n150# a_n417_n150# 0.43fF
C35 a_n129_n150# a_n417_n150# 0.10fF
C36 a_159_n150# a_255_n150# 0.43fF
C37 a_159_n150# a_n465_172# 0.10fF
C38 a_159_n150# a_n225_n150# 0.07fF
C39 a_351_n150# a_255_n150# 0.43fF
C40 a_351_n150# a_n465_172# 0.10fF
C41 a_63_n150# a_255_n150# 0.16fF
C42 a_63_n150# a_n465_172# 0.10fF
C43 a_n225_n150# a_63_n150# 0.10fF
C44 a_n321_n150# a_n465_172# 0.10fF
C45 a_447_n150# w_n647_n360# 0.17fF
C46 a_351_n150# w_n647_n360# 0.10fF
C47 a_255_n150# w_n647_n360# 0.08fF
C48 a_159_n150# w_n647_n360# 0.07fF
C49 a_63_n150# w_n647_n360# 0.04fF
C50 a_n33_n150# w_n647_n360# 0.04fF
C51 a_n129_n150# w_n647_n360# 0.04fF
C52 a_n225_n150# w_n647_n360# 0.07fF
C53 a_n321_n150# w_n647_n360# 0.08fF
C54 a_n417_n150# w_n647_n360# 0.10fF
C55 a_n509_n150# w_n647_n360# 0.17fF
C56 a_n465_172# w_n647_n360# 1.49fF
.ends

.subckt sky130_fd_pr__pfet_01v8_8DL6ZL VSUBS a_n417_n150# a_351_n150# a_255_n150#
+ a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n465_n247# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150# w_n647_n369#
X0 a_63_n150# a_n465_n247# a_n33_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n129_n150# a_n465_n247# a_n225_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n417_n150# a_n465_n247# a_n509_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n33_n150# a_n465_n247# a_n129_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_351_n150# a_n465_n247# a_255_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_255_n150# a_n465_n247# a_159_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n321_n150# a_n465_n247# a_n417_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_159_n150# a_n465_n247# a_63_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n225_n150# a_n465_n247# a_n321_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_447_n150# a_n465_n247# a_351_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n33_n150# a_63_n150# 0.43fF
C1 w_n647_n369# a_n417_n150# 0.07fF
C2 a_159_n150# a_63_n150# 0.43fF
C3 w_n647_n369# a_n33_n150# 0.02fF
C4 w_n647_n369# a_159_n150# 0.04fF
C5 a_n509_n150# a_n417_n150# 0.43fF
C6 a_n225_n150# a_n321_n150# 0.43fF
C7 a_351_n150# a_n465_n247# 0.08fF
C8 a_n225_n150# a_n465_n247# 0.08fF
C9 a_n225_n150# a_n129_n150# 0.43fF
C10 w_n647_n369# a_63_n150# 0.02fF
C11 a_255_n150# a_n129_n150# 0.07fF
C12 a_255_n150# a_n465_n247# 0.08fF
C13 w_n647_n369# a_n509_n150# 0.14fF
C14 a_n33_n150# a_351_n150# 0.07fF
C15 a_159_n150# a_351_n150# 0.16fF
C16 a_n321_n150# a_n465_n247# 0.08fF
C17 a_n129_n150# a_n321_n150# 0.16fF
C18 a_n225_n150# a_n417_n150# 0.16fF
C19 a_159_n150# a_447_n150# 0.10fF
C20 a_n225_n150# a_n33_n150# 0.16fF
C21 a_n225_n150# a_159_n150# 0.07fF
C22 a_n129_n150# a_n465_n247# 0.08fF
C23 a_255_n150# a_n33_n150# 0.10fF
C24 a_255_n150# a_159_n150# 0.43fF
C25 a_63_n150# a_351_n150# 0.10fF
C26 a_63_n150# a_447_n150# 0.07fF
C27 a_n417_n150# a_n321_n150# 0.43fF
C28 w_n647_n369# a_351_n150# 0.07fF
C29 w_n647_n369# a_447_n150# 0.14fF
C30 a_n33_n150# a_n321_n150# 0.10fF
C31 a_n225_n150# a_63_n150# 0.10fF
C32 a_n129_n150# a_n417_n150# 0.10fF
C33 a_n417_n150# a_n465_n247# 0.08fF
C34 w_n647_n369# a_n225_n150# 0.04fF
C35 a_255_n150# a_63_n150# 0.16fF
C36 a_n129_n150# a_n33_n150# 0.43fF
C37 a_n33_n150# a_n465_n247# 0.08fF
C38 w_n647_n369# a_255_n150# 0.05fF
C39 a_n129_n150# a_159_n150# 0.10fF
C40 a_159_n150# a_n465_n247# 0.08fF
C41 a_n225_n150# a_n509_n150# 0.10fF
C42 a_63_n150# a_n321_n150# 0.07fF
C43 w_n647_n369# a_n321_n150# 0.05fF
C44 a_n129_n150# a_63_n150# 0.16fF
C45 a_63_n150# a_n465_n247# 0.08fF
C46 a_n417_n150# a_n33_n150# 0.07fF
C47 w_n647_n369# a_n129_n150# 0.02fF
C48 w_n647_n369# a_n465_n247# 0.47fF
C49 a_n509_n150# a_n321_n150# 0.16fF
C50 a_159_n150# a_n33_n150# 0.16fF
C51 a_351_n150# a_447_n150# 0.43fF
C52 a_n129_n150# a_n509_n150# 0.07fF
C53 a_255_n150# a_351_n150# 0.43fF
C54 a_255_n150# a_447_n150# 0.16fF
C55 a_447_n150# VSUBS 0.03fF
C56 a_351_n150# VSUBS 0.03fF
C57 a_255_n150# VSUBS 0.03fF
C58 a_159_n150# VSUBS 0.03fF
C59 a_63_n150# VSUBS 0.03fF
C60 a_n33_n150# VSUBS 0.03fF
C61 a_n129_n150# VSUBS 0.03fF
C62 a_n225_n150# VSUBS 0.03fF
C63 a_n321_n150# VSUBS 0.03fF
C64 a_n417_n150# VSUBS 0.03fF
C65 a_n509_n150# VSUBS 0.03fF
C66 a_n465_n247# VSUBS 1.07fF
C67 w_n647_n369# VSUBS 4.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EDT3AT a_15_n11# a_n33_n99# w_n211_n221# a_n73_n11#
X0 a_15_n11# a_n33_n99# a_n73_n11# w_n211_n221# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n73_n11# a_n33_n99# 0.02fF
C1 a_15_n11# a_n73_n11# 0.15fF
C2 a_15_n11# a_n33_n99# 0.02fF
C3 a_15_n11# w_n211_n221# 0.09fF
C4 a_n73_n11# w_n211_n221# 0.09fF
C5 a_n33_n99# w_n211_n221# 0.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AQR2CW a_n33_66# a_n78_n106# w_n216_n254# a_20_n106#
X0 a_20_n106# a_n33_66# a_n78_n106# w_n216_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=200000u
C0 a_20_n106# a_n78_n106# 0.21fF
C1 a_20_n106# w_n216_n254# 0.14fF
C2 a_n78_n106# w_n216_n254# 0.14fF
C3 a_n33_66# w_n216_n254# 0.12fF
.ends

.subckt sky130_fd_pr__pfet_01v8_HRYSXS VSUBS a_n33_n211# a_n78_n114# w_n216_n334#
+ a_20_n114#
X0 a_20_n114# a_n33_n211# a_n78_n114# w_n216_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=200000u
C0 w_n216_n334# a_20_n114# 0.20fF
C1 a_n78_n114# w_n216_n334# 0.20fF
C2 a_n78_n114# a_20_n114# 0.42fF
C3 a_20_n114# VSUBS 0.03fF
C4 a_n78_n114# VSUBS 0.03fF
C5 a_n33_n211# VSUBS 0.12fF
C6 w_n216_n334# VSUBS 1.66fF
.ends

.subckt inverter_csvco in vbulkn out vbulkp vdd vss
Xsky130_fd_pr__nfet_01v8_AQR2CW_0 in vss vbulkn out sky130_fd_pr__nfet_01v8_AQR2CW
Xsky130_fd_pr__pfet_01v8_HRYSXS_0 vbulkn in vdd vbulkp out sky130_fd_pr__pfet_01v8_HRYSXS
C0 in vdd 0.01fF
C1 in out 0.11fF
C2 vbulkp vdd 0.04fF
C3 vbulkp out 0.08fF
C4 in vss 0.01fF
C5 vbulkp vbulkn 2.49fF
C6 out vbulkn 0.60fF
C7 vdd vbulkn 0.06fF
C8 in vbulkn 0.54fF
C9 vss vbulkn 0.17fF
.ends

.subckt csvco_branch vctrl in vbp cap_vco_0/t D0 vss out vdd inverter_csvco_0/vss
+ inverter_csvco_0/vdd
Xsky130_fd_pr__nfet_01v8_7H8F5S_0 vctrl inverter_csvco_0/vss inverter_csvco_0/vss
+ vss vss inverter_csvco_0/vss vss vss inverter_csvco_0/vss vss inverter_csvco_0/vss
+ vss vss sky130_fd_pr__nfet_01v8_7H8F5S
Xsky130_fd_pr__pfet_01v8_8DL6ZL_0 vss inverter_csvco_0/vdd inverter_csvco_0/vdd vdd
+ inverter_csvco_0/vdd vdd vdd inverter_csvco_0/vdd vbp vdd inverter_csvco_0/vdd vdd
+ vdd vdd sky130_fd_pr__pfet_01v8_8DL6ZL
Xsky130_fd_pr__nfet_01v8_EDT3AT_0 cap_vco_0/t D0 vss out sky130_fd_pr__nfet_01v8_EDT3AT
Xinverter_csvco_0 in vss out vdd inverter_csvco_0/vdd inverter_csvco_0/vss inverter_csvco
C0 inverter_csvco_0/vdd vdd 1.89fF
C1 out in 0.06fF
C2 in inverter_csvco_0/vss 0.01fF
C3 out cap_vco_0/t 0.70fF
C4 out inverter_csvco_0/vss 0.03fF
C5 in inverter_csvco_0/vdd 0.01fF
C6 vctrl inverter_csvco_0/vss 0.87fF
C7 out inverter_csvco_0/vdd 0.02fF
C8 cap_vco_0/t inverter_csvco_0/vdd 0.10fF
C9 vbp inverter_csvco_0/vdd 0.75fF
C10 out D0 0.09fF
C11 D0 inverter_csvco_0/vss 0.02fF
C12 cap_vco_0/t vdd 0.04fF
C13 vbp vdd 1.21fF
C14 out vss 0.93fF
C15 inverter_csvco_0/vdd vss 0.26fF
C16 in vss 0.69fF
C17 D0 vss -0.67fF
C18 vbp vss 0.13fF
C19 vdd vss 9.58fF
C20 cap_vco_0/t vss 7.22fF
C21 inverter_csvco_0/vss vss 1.79fF
C22 vctrl vss 3.06fF
.ends

.subckt ring_osc vctrl vss vdd csvco_branch_2/vbp csvco_branch_0/inverter_csvco_0/vss
+ D0 csvco_branch_2/cap_vco_0/t out_vco
Xsky130_fd_pr__nfet_01v8_CBAU6Y_0 vss vctrl vss csvco_branch_2/vbp sky130_fd_pr__nfet_01v8_CBAU6Y
Xsky130_fd_pr__pfet_01v8_4757AC_0 vss vdd csvco_branch_2/vbp vdd csvco_branch_2/vbp
+ sky130_fd_pr__pfet_01v8_4757AC
Xcsvco_branch_0 vctrl out_vco csvco_branch_2/vbp csvco_branch_0/cap_vco_0/t D0 vss
+ csvco_branch_1/in vdd csvco_branch_0/inverter_csvco_0/vss csvco_branch_0/inverter_csvco_0/vdd
+ csvco_branch
Xcsvco_branch_2 vctrl csvco_branch_2/in csvco_branch_2/vbp csvco_branch_2/cap_vco_0/t
+ D0 vss out_vco vdd csvco_branch_2/inverter_csvco_0/vss csvco_branch_2/inverter_csvco_0/vdd
+ csvco_branch
Xcsvco_branch_1 vctrl csvco_branch_1/in csvco_branch_2/vbp csvco_branch_1/cap_vco_0/t
+ D0 vss csvco_branch_2/in vdd csvco_branch_1/inverter_csvco_0/vss csvco_branch_1/inverter_csvco_0/vdd
+ csvco_branch
C0 D0 csvco_branch_1/inverter_csvco_0/vss 0.68fF
C1 D0 csvco_branch_0/inverter_csvco_0/vss 0.49fF
C2 csvco_branch_1/in out_vco 0.76fF
C3 csvco_branch_2/in out_vco 0.58fF
C4 D0 csvco_branch_2/inverter_csvco_0/vss 0.68fF
C5 csvco_branch_0/inverter_csvco_0/vss csvco_branch_2/vbp 0.06fF
C6 D0 vctrl 4.41fF
C7 vdd csvco_branch_0/inverter_csvco_0/vdd 0.13fF
C8 csvco_branch_1/inverter_csvco_0/vdd vdd 0.19fF
C9 vdd csvco_branch_2/inverter_csvco_0/vdd 0.10fF
C10 vctrl csvco_branch_2/vbp 0.06fF
C11 csvco_branch_2/vbp csvco_branch_0/inverter_csvco_0/vdd 0.06fF
C12 out_vco csvco_branch_1/cap_vco_0/t 0.03fF
C13 out_vco csvco_branch_0/cap_vco_0/t 0.03fF
C14 vdd csvco_branch_2/vbp 1.49fF
C15 csvco_branch_2/in vss 1.60fF
C16 csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C17 csvco_branch_1/cap_vco_0/t vss 7.10fF
C18 csvco_branch_1/inverter_csvco_0/vss vss 0.72fF
C19 csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C20 csvco_branch_2/cap_vco_0/t vss 7.10fF
C21 csvco_branch_2/inverter_csvco_0/vss vss 0.62fF
C22 csvco_branch_1/in vss 1.58fF
C23 csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C24 out_vco vss 0.67fF
C25 D0 vss -1.55fF
C26 vdd vss 31.40fF
C27 csvco_branch_0/cap_vco_0/t vss 7.10fF
C28 csvco_branch_0/inverter_csvco_0/vss vss 0.66fF
C29 vctrl vss 11.02fF
C30 csvco_branch_2/vbp vss 0.77fF
.ends

.subckt ring_osc_buffer vss in_vco vdd o1 out_div out_pad
Xinverter_min_x4_0 o1 vss out_div vdd inverter_min_x4
Xinverter_min_x4_1 out_div vss out_pad vdd inverter_min_x4
Xinverter_min_x2_0 in_vco o1 vss vdd inverter_min_x2
C0 vdd out_pad 0.10fF
C1 o1 out_div 0.11fF
C2 out_pad out_div 0.15fF
C3 vdd out_div 0.17fF
C4 vdd o1 0.09fF
C5 vdd vss 14.54fF
C6 in_vco vss 0.83fF
C7 out_pad vss 0.70fF
C8 out_div vss 3.00fF
C9 o1 vss 2.72fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AZESM8 a_n63_n151# a_n33_n125# a_n255_n151# a_33_n151#
+ a_n225_n125# a_63_n125# a_n129_n125# a_n159_n151# w_n455_n335# a_225_n151# a_255_n125#
+ a_129_n151# a_159_n125# a_n317_n125#
X0 a_159_n125# a_129_n151# a_63_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n225_n125# a_n255_n151# a_n317_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_63_n125# a_33_n151# a_n33_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_n129_n125# a_n159_n151# a_n225_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n33_n125# a_n63_n151# a_n129_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_255_n125# a_225_n151# a_159_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n63_n151# a_n159_n151# 0.02fF
C1 a_n63_n151# a_33_n151# 0.02fF
C2 a_225_n151# a_129_n151# 0.02fF
C3 a_159_n125# a_255_n125# 0.36fF
C4 a_n129_n125# a_159_n125# 0.08fF
C5 a_n159_n151# a_n255_n151# 0.02fF
C6 a_159_n125# a_n33_n125# 0.13fF
C7 a_n129_n125# a_n317_n125# 0.13fF
C8 a_63_n125# a_255_n125# 0.13fF
C9 a_n317_n125# a_n33_n125# 0.08fF
C10 a_n129_n125# a_63_n125# 0.13fF
C11 a_n129_n125# a_n225_n125# 0.36fF
C12 a_63_n125# a_n33_n125# 0.36fF
C13 a_n225_n125# a_n33_n125# 0.13fF
C14 a_159_n125# a_63_n125# 0.36fF
C15 a_159_n125# a_n225_n125# 0.06fF
C16 a_129_n151# a_33_n151# 0.02fF
C17 a_n317_n125# a_63_n125# 0.06fF
C18 a_n317_n125# a_n225_n125# 0.36fF
C19 a_n129_n125# a_255_n125# 0.06fF
C20 a_255_n125# a_n33_n125# 0.08fF
C21 a_63_n125# a_n225_n125# 0.08fF
C22 a_n129_n125# a_n33_n125# 0.36fF
C23 a_255_n125# w_n455_n335# 0.14fF
C24 a_159_n125# w_n455_n335# 0.08fF
C25 a_63_n125# w_n455_n335# 0.07fF
C26 a_n33_n125# w_n455_n335# 0.08fF
C27 a_n129_n125# w_n455_n335# 0.07fF
C28 a_n225_n125# w_n455_n335# 0.08fF
C29 a_n317_n125# w_n455_n335# 0.14fF
C30 a_225_n151# w_n455_n335# 0.05fF
C31 a_129_n151# w_n455_n335# 0.05fF
C32 a_33_n151# w_n455_n335# 0.05fF
C33 a_n63_n151# w_n455_n335# 0.05fF
C34 a_n159_n151# w_n455_n335# 0.05fF
C35 a_n255_n151# w_n455_n335# 0.05fF
.ends

.subckt sky130_fd_pr__pfet_01v8_XJXT7S VSUBS a_n33_n125# a_n255_n154# a_33_n154# a_n225_n125#
+ a_n159_n154# a_63_n125# a_n129_n125# a_225_n154# a_129_n154# a_255_n125# a_159_n125#
+ a_n317_n125# w_n455_n344# a_n63_n154#
X0 a_n129_n125# a_n159_n154# a_n225_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n33_n125# a_n63_n154# a_n129_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_255_n125# a_225_n154# a_159_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_159_n125# a_129_n154# a_63_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n225_n125# a_n255_n154# a_n317_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_63_n125# a_33_n154# a_n33_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_63_n125# a_255_n125# 0.13fF
C1 a_63_n125# a_n33_n125# 0.36fF
C2 a_63_n125# a_n129_n125# 0.13fF
C3 a_n225_n125# a_n33_n125# 0.13fF
C4 a_n129_n125# a_n225_n125# 0.36fF
C5 a_63_n125# a_n225_n125# 0.08fF
C6 w_n455_n344# a_159_n125# 0.06fF
C7 a_n63_n154# a_33_n154# 0.02fF
C8 a_n159_n154# a_n255_n154# 0.02fF
C9 a_n317_n125# a_n33_n125# 0.08fF
C10 a_129_n154# a_225_n154# 0.02fF
C11 a_n317_n125# a_n129_n125# 0.13fF
C12 w_n455_n344# a_255_n125# 0.11fF
C13 w_n455_n344# a_n33_n125# 0.05fF
C14 w_n455_n344# a_n129_n125# 0.04fF
C15 a_n317_n125# a_63_n125# 0.06fF
C16 w_n455_n344# a_63_n125# 0.04fF
C17 a_n317_n125# a_n225_n125# 0.36fF
C18 w_n455_n344# a_n225_n125# 0.06fF
C19 a_n63_n154# a_n159_n154# 0.02fF
C20 a_159_n125# a_255_n125# 0.36fF
C21 a_159_n125# a_n33_n125# 0.13fF
C22 a_159_n125# a_n129_n125# 0.08fF
C23 a_n317_n125# w_n455_n344# 0.11fF
C24 a_63_n125# a_159_n125# 0.36fF
C25 a_129_n154# a_33_n154# 0.02fF
C26 a_159_n125# a_n225_n125# 0.06fF
C27 a_n33_n125# a_255_n125# 0.08fF
C28 a_n129_n125# a_255_n125# 0.06fF
C29 a_n129_n125# a_n33_n125# 0.36fF
C30 a_255_n125# VSUBS 0.03fF
C31 a_159_n125# VSUBS 0.03fF
C32 a_63_n125# VSUBS 0.03fF
C33 a_n33_n125# VSUBS 0.03fF
C34 a_n129_n125# VSUBS 0.03fF
C35 a_n225_n125# VSUBS 0.03fF
C36 a_n317_n125# VSUBS 0.03fF
C37 a_225_n154# VSUBS 0.05fF
C38 a_129_n154# VSUBS 0.05fF
C39 a_33_n154# VSUBS 0.05fF
C40 a_n63_n154# VSUBS 0.05fF
C41 a_n159_n154# VSUBS 0.05fF
C42 a_n255_n154# VSUBS 0.05fF
C43 w_n455_n344# VSUBS 2.96fF
.ends

.subckt inverter_cp_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_AZESM8_0 in vss in in vss out out in vss in out in vss out
+ sky130_fd_pr__nfet_01v8_AZESM8
Xsky130_fd_pr__pfet_01v8_XJXT7S_0 vss vdd in in vdd in out out in in out vdd out vdd
+ in sky130_fd_pr__pfet_01v8_XJXT7S
C0 out in 0.85fF
C1 vdd in 0.04fF
C2 vdd out 0.29fF
C3 vdd vss 5.90fF
C4 out vss 1.30fF
C5 in vss 1.82fF
.ends

.subckt pfd_cp_interface vss vdd inverter_cp_x1_0/out inverter_cp_x1_2/in Down QA
+ QB nDown Up nUp
Xinverter_cp_x2_0 nDown Down vss vdd inverter_cp_x2
Xinverter_cp_x2_1 Up nUp vss vdd inverter_cp_x2
Xtrans_gate_0 nDown vss inverter_cp_x1_0/out vdd trans_gate
Xinverter_cp_x1_0 inverter_cp_x1_0/out QB vss vdd inverter_cp_x1
Xinverter_cp_x1_1 inverter_cp_x1_2/in QA vss vdd inverter_cp_x1
Xinverter_cp_x1_2 Up inverter_cp_x1_2/in vss vdd inverter_cp_x1
C0 vdd nUp 0.14fF
C1 nUp Up 0.20fF
C2 vdd QA 0.02fF
C3 vdd inverter_cp_x1_2/in 0.42fF
C4 vdd QB 0.02fF
C5 inverter_cp_x1_2/in Up 0.12fF
C6 Down inverter_cp_x1_0/out 0.12fF
C7 vdd inverter_cp_x1_0/out 0.18fF
C8 vdd Up 0.60fF
C9 nDown Down 0.23fF
C10 vdd nDown 0.80fF
C11 nDown inverter_cp_x1_0/out 0.11fF
C12 inverter_cp_x1_2/in vss 2.01fF
C13 QA vss 1.09fF
C14 inverter_cp_x1_0/out vss 1.72fF
C15 QB vss 1.09fF
C16 vdd vss 28.20fF
C17 nUp vss 1.32fF
C18 Up vss 2.53fF
C19 Down vss 1.17fF
C20 nDown vss 2.77fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4F35BC VSUBS a_n129_n90# w_n359_n309# a_n63_n116#
+ a_n159_n207# a_63_n90# a_n33_n90# a_n221_n90# a_159_n90#
X0 a_159_n90# a_n63_n116# a_63_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n129_n90# a_n159_n207# a_n221_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X2 a_63_n90# a_n159_n207# a_n33_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3 a_n33_n90# a_n63_n116# a_n129_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_n129_n90# a_n221_n90# 0.26fF
C1 a_63_n90# a_n221_n90# 0.06fF
C2 a_n129_n90# a_159_n90# 0.06fF
C3 a_n33_n90# w_n359_n309# 0.05fF
C4 a_63_n90# a_159_n90# 0.26fF
C5 w_n359_n309# a_n221_n90# 0.09fF
C6 a_n33_n90# a_n221_n90# 0.09fF
C7 a_159_n90# w_n359_n309# 0.09fF
C8 a_159_n90# a_n33_n90# 0.09fF
C9 a_63_n90# a_n129_n90# 0.09fF
C10 a_n63_n116# a_n159_n207# 0.12fF
C11 a_159_n90# a_n221_n90# 0.04fF
C12 a_n129_n90# w_n359_n309# 0.06fF
C13 a_n129_n90# a_n33_n90# 0.26fF
C14 a_63_n90# w_n359_n309# 0.06fF
C15 a_63_n90# a_n33_n90# 0.26fF
C16 a_159_n90# VSUBS 0.03fF
C17 a_63_n90# VSUBS 0.03fF
C18 a_n33_n90# VSUBS 0.03fF
C19 a_n129_n90# VSUBS 0.03fF
C20 a_n221_n90# VSUBS 0.03fF
C21 a_n159_n207# VSUBS 0.30fF
C22 a_n63_n116# VSUBS 0.37fF
C23 w_n359_n309# VSUBS 2.23fF
.ends

.subckt sky130_fd_pr__nfet_01v8_C3YG4M a_n33_n45# a_33_n71# a_n129_71# w_n263_n255#
+ a_n125_n45# a_63_n45#
X0 a_63_n45# a_33_n71# a_n33_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n129_71# a_n125_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_n129_71# a_33_n71# 0.04fF
C1 a_63_n45# a_n125_n45# 0.05fF
C2 a_63_n45# a_n33_n45# 0.13fF
C3 a_n125_n45# a_n33_n45# 0.13fF
C4 a_63_n45# w_n263_n255# 0.04fF
C5 a_n33_n45# w_n263_n255# 0.04fF
C6 a_n125_n45# w_n263_n255# 0.04fF
C7 a_33_n71# w_n263_n255# 0.11fF
C8 a_n129_71# w_n263_n255# 0.14fF
.ends

.subckt nor_pfd vdd sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss A B
Xsky130_fd_pr__pfet_01v8_4F35BC_0 vss sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vdd B A sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out vdd vdd sky130_fd_pr__pfet_01v8_4F35BC
Xsky130_fd_pr__nfet_01v8_C3YG4M_0 out B A vss vss vss sky130_fd_pr__nfet_01v8_C3YG4M
C0 out B 0.40fF
C1 A B 0.24fF
C2 vdd out 0.11fF
C3 A out 0.06fF
C4 vdd sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.02fF
C5 vdd A 0.09fF
C6 sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out 0.08fF
C7 vdd sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.02fF
C8 sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C9 out vss 0.45fF
C10 sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C11 A vss 0.83fF
C12 B vss 1.09fF
C13 vdd vss 3.79fF
.ends

.subckt dff_pfd vss vdd nor_pfd_2/A Q CLK nor_pfd_3/A Reset nor_pfd_2/B
Xnor_pfd_0 vdd nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_2/A nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss CLK Q nor_pfd
Xnor_pfd_1 vdd nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# Q nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss nor_pfd_2/A nor_pfd_3/A nor_pfd
Xnor_pfd_2 vdd nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_3/A nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss nor_pfd_2/A nor_pfd_2/B nor_pfd
Xnor_pfd_3 vdd nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_2/B nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss nor_pfd_3/A Reset nor_pfd
C0 Q nor_pfd_3/A 0.98fF
C1 vdd nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.06fF
C2 Q CLK 0.04fF
C3 vdd nor_pfd_2/A -0.01fF
C4 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vdd 0.06fF
C5 vdd nor_pfd_2/B 0.02fF
C6 vdd nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.06fF
C7 Q nor_pfd_2/A 1.38fF
C8 Q nor_pfd_2/B 2.22fF
C9 Q Reset 0.14fF
C10 vdd nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.06fF
C11 vdd nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.06fF
C12 nor_pfd_3/A nor_pfd_2/A 0.38fF
C13 nor_pfd_3/A nor_pfd_2/B 0.58fF
C14 vdd Q 0.08fF
C15 nor_pfd_3/A Reset 0.12fF
C16 nor_pfd_2/A nor_pfd_2/B 0.05fF
C17 Reset nor_pfd_2/B 0.43fF
C18 vdd nor_pfd_3/A 0.09fF
C19 vdd nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.06fF
C20 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C21 nor_pfd_2/B vss 1.42fF
C22 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C23 nor_pfd_3/A vss 3.16fF
C24 Reset vss 1.48fF
C25 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C26 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C27 nor_pfd_2/A vss 2.56fF
C28 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C29 Q vss 2.77fF
C30 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C31 vdd vss 16.42fF
C32 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C33 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C34 CLK vss 0.95fF
.ends

.subckt sky130_fd_pr__nfet_01v8_ZCYAJJ w_n359_n255# a_n33_n45# a_n159_n173# a_n221_n45#
+ a_159_n45# a_n63_n71# a_n129_n45# a_63_n45#
X0 a_63_n45# a_n159_n173# a_n33_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n63_n71# a_n129_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X2 a_159_n45# a_n63_n71# a_63_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X3 a_n129_n45# a_n159_n173# a_n221_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_63_n45# a_n33_n45# 0.13fF
C1 a_159_n45# a_n221_n45# 0.02fF
C2 a_159_n45# a_63_n45# 0.13fF
C3 a_159_n45# a_n33_n45# 0.05fF
C4 a_n221_n45# a_n129_n45# 0.13fF
C5 a_63_n45# a_n129_n45# 0.05fF
C6 a_n159_n173# a_n63_n71# 0.10fF
C7 a_n129_n45# a_n33_n45# 0.13fF
C8 a_63_n45# a_n221_n45# 0.03fF
C9 a_159_n45# a_n129_n45# 0.03fF
C10 a_n221_n45# a_n33_n45# 0.05fF
C11 a_159_n45# w_n359_n255# 0.04fF
C12 a_63_n45# w_n359_n255# 0.05fF
C13 a_n33_n45# w_n359_n255# 0.05fF
C14 a_n129_n45# w_n359_n255# 0.05fF
C15 a_n221_n45# w_n359_n255# 0.08fF
C16 a_n159_n173# w_n359_n255# 0.31fF
C17 a_n63_n71# w_n359_n255# 0.31fF
.ends

.subckt sky130_fd_pr__pfet_01v8_7T83YG VSUBS a_n125_n90# a_63_n90# a_33_n187# a_n99_n187#
+ a_n33_n90# w_n263_n309#
X0 a_63_n90# a_33_n187# a_n33_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n33_n90# a_n99_n187# a_n125_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_n125_n90# a_n33_n90# 0.26fF
C1 a_n99_n187# a_33_n187# 0.04fF
C2 a_n125_n90# a_63_n90# 0.09fF
C3 a_n33_n90# a_63_n90# 0.26fF
C4 a_63_n90# VSUBS 0.03fF
C5 a_n33_n90# VSUBS 0.03fF
C6 a_n125_n90# VSUBS 0.03fF
C7 a_33_n187# VSUBS 0.12fF
C8 a_n99_n187# VSUBS 0.12fF
C9 w_n263_n309# VSUBS 1.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_ZXAV3F a_n73_n45# a_n33_67# a_15_n45# w_n211_n255#
X0 a_15_n45# a_n33_67# a_n73_n45# w_n211_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_n73_n45# a_15_n45# 0.16fF
C1 a_15_n45# w_n211_n255# 0.08fF
C2 a_n73_n45# w_n211_n255# 0.06fF
C3 a_n33_67# w_n211_n255# 0.10fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4F7GBC VSUBS a_n51_n187# a_n73_n90# a_15_n90# w_n211_n309#
X0 a_15_n90# a_n51_n187# a_n73_n90# w_n211_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_15_n90# w_n211_n309# 0.09fF
C1 a_n73_n90# w_n211_n309# 0.04fF
C2 a_15_n90# a_n73_n90# 0.31fF
C3 a_15_n90# VSUBS 0.03fF
C4 a_n73_n90# VSUBS 0.03fF
C5 a_n51_n187# VSUBS 0.12fF
C6 w_n211_n309# VSUBS 1.24fF
.ends

.subckt and_pfd a_656_410# out vss vdd A B
Xsky130_fd_pr__nfet_01v8_ZCYAJJ_0 vss a_656_410# A vss vss B sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45#
+ sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# sky130_fd_pr__nfet_01v8_ZCYAJJ
Xsky130_fd_pr__pfet_01v8_7T83YG_0 vss vdd vdd B A a_656_410# vdd sky130_fd_pr__pfet_01v8_7T83YG
Xsky130_fd_pr__nfet_01v8_ZXAV3F_0 vss a_656_410# out vss sky130_fd_pr__nfet_01v8_ZXAV3F
Xsky130_fd_pr__pfet_01v8_4F7GBC_0 vss a_656_410# vdd out vdd sky130_fd_pr__pfet_01v8_4F7GBC
C0 vdd out 0.10fF
C1 A a_656_410# 0.04fF
C2 a_656_410# out 0.20fF
C3 A B 0.33fF
C4 a_656_410# sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# 0.07fF
C5 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# B 0.02fF
C6 out sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# 0.03fF
C7 vdd a_656_410# 0.20fF
C8 a_656_410# B 0.30fF
C9 A vdd 0.05fF
C10 vdd vss 4.85fF
C11 out vss 0.47fF
C12 a_656_410# vss 1.00fF
C13 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.13fF
C14 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.10fF
C15 A vss 0.85fF
C16 B vss 0.95fF
.ends

.subckt PFD vss vdd Reset Down Up A B
Xdff_pfd_0 vss vdd dff_pfd_0/nor_pfd_2/A Up A dff_pfd_0/nor_pfd_3/A Reset dff_pfd_0/nor_pfd_2/B
+ dff_pfd
Xdff_pfd_1 vss vdd dff_pfd_1/nor_pfd_2/A Down B dff_pfd_1/nor_pfd_3/A Reset dff_pfd_1/nor_pfd_2/B
+ dff_pfd
Xand_pfd_0 and_pfd_0/a_656_410# Reset vss vdd Up Down and_pfd
C0 vdd dff_pfd_0/nor_pfd_2/A 0.13fF
C1 dff_pfd_0/nor_pfd_3/A vdd 0.08fF
C2 Up vdd 1.62fF
C3 Up Down 0.06fF
C4 dff_pfd_1/nor_pfd_3/A vdd 0.08fF
C5 dff_pfd_1/nor_pfd_2/B vdd 0.04fF
C6 dff_pfd_1/nor_pfd_2/A vdd 0.13fF
C7 dff_pfd_0/nor_pfd_2/B vdd 0.11fF
C8 Down vdd 0.08fF
C9 Reset vdd 0.02fF
C10 and_pfd_0/a_656_410# vss 0.99fF
C11 and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C12 and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.05fF
C13 dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C14 dff_pfd_1/nor_pfd_2/B vss 1.51fF
C15 dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C16 dff_pfd_1/nor_pfd_3/A vss 3.14fF
C17 dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C18 dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C19 dff_pfd_1/nor_pfd_2/A vss 2.56fF
C20 dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C21 Down vss 3.74fF
C22 dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C23 vdd vss 44.73fF
C24 dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C25 dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C26 B vss 1.07fF
C27 dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C28 dff_pfd_0/nor_pfd_2/B vss 1.40fF
C29 dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C30 dff_pfd_0/nor_pfd_3/A vss 3.14fF
C31 Reset vss 3.85fF
C32 dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C33 dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C34 dff_pfd_0/nor_pfd_2/A vss 2.56fF
C35 dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C36 Up vss 3.18fF
C37 dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C38 dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C39 dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C40 A vss 1.07fF
.ends


* Top level circuit top_pll_v3

Xcharge_pump_0 nswitch vss vdd nUp Down charge_pump_0/w_2544_775# vco_vctrl pswitch
+ iref_cp nDown biasp Up vss charge_pump
Xloop_filter_v2_0 lf_vc lf_D0 vco_vctrl vss loop_filter_v2
Xdiv_by_2_0 vdd vss n_out_div_2 out_by_2 n_out_by_2 out_buffer_div_2 n_out_buffer_div_2
+ out_to_div out_div_2 div_by_2
Xfreq_div_0 clk_0 vss n_clk_0 vdd freq_div_0/prescaler_23_0/Q2 s_0 s_1_n s_1 freq_div_0/prescaler_23_0/nCLK_23
+ MC clk_d freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# s_0_n clk_pre
+ freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/D
+ freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/nD clk_1 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280#
+ clk_out_mux21 n_clk_1 out_div freq_div_0/div_by_5_0/Q1 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D
+ freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD
+ clk_2_f out_by_2 n_out_by_2 clk_5 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/D
+ freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/nD freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D
+ freq_div
Xbuffer_salida_0 buffer_salida_0/a_678_n100# out_to_pad vdd out_to_buffer vss buffer_salida
Xring_osc_0 vco_vctrl vss vdd ring_osc_0/csvco_branch_2/vbp ring_osc_0/csvco_branch_0/inverter_csvco_0/vss
+ vco_D0 ring_osc_0/csvco_branch_2/cap_vco_0/t vco_out ring_osc
Xring_osc_buffer_0 vss vco_out vdd out_first_buffer out_to_div out_to_buffer ring_osc_buffer
Xpfd_cp_interface_0 vss vdd pfd_cp_interface_0/inverter_cp_x1_0/out pfd_cp_interface_0/inverter_cp_x1_2/in
+ Down QA QB nDown Up nUp pfd_cp_interface
XPFD_0 vss vdd pfd_reset QB QA in_ref out_div PFD
C0 vco_vctrl freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/D 0.53fF
C1 biasp nUp -0.16fF
C2 iref_cp Down 0.09fF
C3 vco_vctrl freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/D 0.09fF
C4 vco_vctrl freq_div_0/prescaler_23_0/Q2 0.06fF
C5 clk_d out_div 0.60fF
C6 vco_vctrl vdd 0.58fF
C7 vco_vctrl freq_div_0/div_by_5_0/Q1 0.10fF
C8 ring_osc_0/csvco_branch_2/vbp vco_vctrl 0.26fF
C9 vdd nUp 0.05fF
C10 vco_vctrl n_clk_1 0.23fF
C11 MC vco_vctrl 0.33fF
C12 charge_pump_0/w_2544_775# nDown 0.05fF
C13 Down nDown 2.55fF
C14 QA vdd -0.04fF
C15 vco_vctrl s_0_n 0.34fF
C16 vco_vctrl freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD 0.15fF
C17 nswitch nDown 0.76fF
C18 vco_vctrl clk_0 -0.26fF
C19 ring_osc_0/csvco_branch_2/vbp vdd 0.03fF
C20 pswitch Up 1.98fF
C21 vco_vctrl freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D -0.42fF
C22 nUp Up 2.72fF
C23 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/nD vco_vctrl 0.09fF
C24 out_to_buffer vdd 0.07fF
C25 vco_vctrl freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD -0.42fF
C26 vco_vctrl s_0 0.45fF
C27 biasp Down 1.24fF
C28 n_out_by_2 s_0_n 0.14fF
C29 ring_osc_0/csvco_branch_2/cap_vco_0/t vdd 0.02fF
C30 biasp Up 0.26fF
C31 MC lf_vc 0.20fF
C32 out_by_2 n_out_by_2 0.27fF
C33 clk_0 vdd 0.13fF
C34 vdd Up 0.28fF
C35 pfd_cp_interface_0/inverter_cp_x1_2/in vdd 0.01fF
C36 vdd buffer_salida_0/a_678_n100# 0.24fF
C37 n_out_by_2 s_0 0.14fF
C38 charge_pump_0/w_2544_775# Down -0.23fF
C39 vco_vctrl clk_1 -0.04fF
C40 out_to_buffer buffer_salida_0/a_678_n100# 0.21fF
C41 vco_vctrl freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D 0.65fF
C42 nswitch Down 0.54fF
C43 out_to_buffer out_to_div 0.13fF
C44 s_1 out_div 0.37fF
C45 pswitch nDown 0.53fF
C46 nDown nUp -0.09fF
C47 n_out_by_2 clk_1 -0.10fF
C48 vco_D0 vdd 0.03fF
C49 vco_vctrl freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# 0.82fF
C50 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# vco_vctrl 0.17fF
C51 pswitch nUp 0.93fF
C52 ring_osc_0/csvco_branch_2/cap_vco_0/t out_first_buffer 0.03fF
C53 vco_vctrl ring_osc_0/csvco_branch_0/inverter_csvco_0/vss 0.04fF
C54 vco_vctrl freq_div_0/prescaler_23_0/nCLK_23 0.06fF
C55 biasp nDown 0.26fF
C56 vco_vctrl freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# 0.34fF
C57 out_to_div s_0 0.94fF
C58 s_1_n out_div 0.09fF
C59 vdd nDown 0.22fF
C60 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/nD vco_vctrl 1.23fF
C61 PFD_0/and_pfd_0/a_656_410# vss 0.96fF
C62 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C63 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.07fF
C64 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C65 PFD_0/dff_pfd_1/nor_pfd_2/B vss 1.40fF
C66 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C67 PFD_0/dff_pfd_1/nor_pfd_3/A vss 3.14fF
C68 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C69 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C70 PFD_0/dff_pfd_1/nor_pfd_2/A vss 2.55fF
C71 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C72 QB vss 3.15fF
C73 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C74 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C75 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C76 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C77 PFD_0/dff_pfd_0/nor_pfd_2/B vss 1.40fF
C78 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C79 PFD_0/dff_pfd_0/nor_pfd_3/A vss 3.14fF
C80 pfd_reset vss 1.87fF
C81 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C82 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C83 PFD_0/dff_pfd_0/nor_pfd_2/A vss 2.55fF
C84 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C85 QA vss 3.49fF
C86 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C87 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C88 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C89 in_ref vss 0.84fF
C90 pfd_cp_interface_0/inverter_cp_x1_2/in vss 1.85fF
C91 pfd_cp_interface_0/inverter_cp_x1_0/out vss 1.66fF
C92 nUp vss 0.12fF
C93 Up vss -4.26fF
C94 Down vss 1.89fF
C95 nDown vss 2.59fF
C96 out_to_buffer vss 1.92fF
C97 out_to_div vss 8.72fF
C98 out_first_buffer vss 2.15fF
C99 ring_osc_0/csvco_branch_2/in vss 1.60fF
C100 ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C101 ring_osc_0/csvco_branch_1/cap_vco_0/t vss 7.10fF
C102 ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vss 0.52fF
C103 ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C104 ring_osc_0/csvco_branch_2/cap_vco_0/t vss 7.10fF
C105 ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vss 0.52fF
C106 ring_osc_0/csvco_branch_1/in vss 1.58fF
C107 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C108 vco_out vss 1.65fF
C109 vco_D0 vss -4.72fF
C110 ring_osc_0/csvco_branch_0/cap_vco_0/t vss 7.10fF
C111 ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vss 0.52fF
C112 ring_osc_0/csvco_branch_2/vbp vss 0.38fF
C113 out_to_pad vss 7.15fF
C114 buffer_salida_0/a_3996_n100# vss 48.29fF
C115 buffer_salida_0/a_678_n100# vss 13.38fF
C116 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_1/a_63_368# vss 0.37fF
C117 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C118 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_0/X vss 0.49fF
C119 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C120 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C121 freq_div_0/prescaler_23_0/Q2_d vss -0.69fF
C122 freq_div_0/prescaler_23_0/DFlipFlop_2/nQ vss 0.48fF
C123 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C124 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C125 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C126 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C127 freq_div_0/prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C128 freq_div_0/prescaler_23_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C129 freq_div_0/prescaler_23_0/Q2 vss 0.55fF
C130 freq_div_0/prescaler_23_0/DFlipFlop_2/latch_diff_0/nD vss 0.94fF
C131 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C132 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C133 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C134 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C135 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C136 freq_div_0/prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C137 freq_div_0/prescaler_23_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C138 freq_div_0/prescaler_23_0/DFlipFlop_1/D vss 1.90fF
C139 freq_div_0/prescaler_23_0/DFlipFlop_1/latch_diff_0/nD vss 0.94fF
C140 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C141 n_clk_0 vss -6.63fF
C142 freq_div_0/prescaler_23_0/Q1 vss 0.07fF
C143 freq_div_0/prescaler_23_0/DFlipFlop_0/nQ vss 0.48fF
C144 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C145 clk_0 vss -0.36fF
C146 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C147 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C148 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C149 freq_div_0/prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C150 freq_div_0/prescaler_23_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C151 freq_div_0/prescaler_23_0/nCLK_23 vss -1.02fF
C152 freq_div_0/prescaler_23_0/DFlipFlop_0/latch_diff_0/nD vss 0.94fF
C153 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__or2_1_1/X vss -1.01fF
C154 MC vss -1.42fF
C155 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_304_74# vss 0.36fF
C156 freq_div_0/prescaler_23_0/sky130_fd_sc_hs__mux2_1_0/a_27_112# vss 0.65fF
C157 n_out_by_2 vss 4.53fF
C158 out_by_2 vss 4.18fF
C159 s_0_n vss -3.95fF
C160 s_0 vss 5.61fF
C161 freq_div_0/div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C162 freq_div_0/div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.38fF
C163 freq_div_0/div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C164 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.57fF
C165 freq_div_0/div_by_5_0/Q1_shift vss -0.36fF
C166 freq_div_0/div_by_5_0/DFlipFlop_3/nQ vss 0.48fF
C167 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C168 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_1/D vss -1.73fF
C169 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C170 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_0/D vss 0.96fF
C171 freq_div_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C172 freq_div_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C173 freq_div_0/div_by_5_0/Q1 vss 4.35fF
C174 freq_div_0/div_by_5_0/DFlipFlop_3/latch_diff_0/nD vss 0.94fF
C175 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C176 freq_div_0/div_by_5_0/Q0 vss 0.29fF
C177 freq_div_0/div_by_5_0/nQ0 vss 0.99fF
C178 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C179 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C180 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C181 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C182 freq_div_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C183 freq_div_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C184 freq_div_0/div_by_5_0/DFlipFlop_1/D vss 3.64fF
C185 freq_div_0/div_by_5_0/DFlipFlop_1/latch_diff_0/nD vss 0.94fF
C186 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C187 freq_div_0/div_by_5_0/DFlipFlop_2/nQ vss 0.48fF
C188 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C189 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C190 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C191 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C192 freq_div_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C193 freq_div_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C194 freq_div_0/div_by_5_0/DFlipFlop_2/D vss 3.13fF
C195 freq_div_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD vss 0.94fF
C196 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C197 n_clk_1 vss -0.57fF
C198 freq_div_0/div_by_5_0/DFlipFlop_0/Q vss -0.94fF
C199 freq_div_0/div_by_5_0/nQ2 vss 1.38fF
C200 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C201 clk_1 vss -2.22fF
C202 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C203 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C204 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C205 freq_div_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C206 freq_div_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C207 freq_div_0/div_by_5_0/DFlipFlop_0/D vss 3.96fF
C208 vdd vss 573.83fF
C209 freq_div_0/div_by_5_0/DFlipFlop_0/latch_diff_0/nD vss 0.94fF
C210 freq_div_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C211 freq_div_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.40fF
C212 out_div vss 3.34fF
C213 clk_d vss 1.26fF
C214 s_1_n vss -2.01fF
C215 s_1 vss 1.77fF
C216 freq_div_0/inverter_min_x4_0/in vss 2.71fF
C217 clk_5 vss -0.23fF
C218 clk_out_mux21 vss 3.65fF
C219 clk_pre vss 1.67fF
C220 clk_2_f vss 3.29fF
C221 freq_div_0/div_by_2_0/o1 vss 2.08fF
C222 freq_div_0/div_by_2_0/nCLK_2 vss 1.04fF
C223 freq_div_0/div_by_2_0/o2 vss 2.08fF
C224 freq_div_0/div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C225 freq_div_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C226 freq_div_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C227 freq_div_0/div_by_2_0/DFlipFlop_0/nCLK vss 0.82fF
C228 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C229 freq_div_0/div_by_2_0/out_div vss -0.82fF
C230 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C231 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C232 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C233 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C234 freq_div_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C235 freq_div_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C236 freq_div_0/div_by_2_0/nout_div vss 2.62fF
C237 freq_div_0/div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 0.94fF
C238 out_buffer_div_2 vss 1.57fF
C239 n_out_buffer_div_2 vss 1.57fF
C240 div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C241 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C242 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C243 div_by_2_0/DFlipFlop_0/nCLK vss 0.82fF
C244 div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C245 out_div_2 vss -0.70fF
C246 div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C247 div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C248 div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C249 div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C250 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C251 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.56fF
C252 n_out_div_2 vss 2.11fF
C253 div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 0.94fF
C254 lf_vc vss -60.88fF
C255 loop_filter_v2_0/res_loop_filter_2/out vss 7.90fF
C256 lf_D0 vss 0.01fF
C257 loop_filter_v2_0/cap3_loop_filter_0/in vss -12.03fF
C258 nswitch vss 4.61fF
C259 biasp vss 5.46fF
C260 iref_cp vss 2.44fF
C261 vco_vctrl vss -30.43fF
C262 pswitch vss 2.72fF
.end

