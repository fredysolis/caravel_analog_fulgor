magic
tech sky130A
magscale 1 2
timestamp 1623892191
<< error_p >>
rect -8209 8140 -7989 13200
rect -13288 8000 -7989 8140
rect -7969 8140 -7749 13200
rect -2890 8140 -2670 13200
rect -7969 8000 -2670 8140
rect -2650 8140 -2430 13200
rect 2429 8140 2649 13200
rect -2650 8000 2649 8140
rect 2669 8140 2889 13200
rect 7748 8140 7968 13200
rect 2669 8000 7968 8140
rect 7988 8140 8208 13200
rect 7988 8000 13287 8140
rect -13288 7760 -7989 7900
rect -8209 2840 -7989 7760
rect -13288 2700 -7989 2840
rect -7969 7760 -2670 7900
rect -7969 2840 -7749 7760
rect -2890 2840 -2670 7760
rect -7969 2700 -2670 2840
rect -2650 7760 2649 7900
rect -2650 2840 -2430 7760
rect 2429 2840 2649 7760
rect -2650 2700 2649 2840
rect 2669 7760 7968 7900
rect 2669 2840 2889 7760
rect 7748 2840 7968 7760
rect 2669 2700 7968 2840
rect 7988 7760 13287 7900
rect 7988 2840 8208 7760
rect 7988 2700 13287 2840
rect -13288 2460 -7989 2600
rect -8209 -2460 -7989 2460
rect -13288 -2600 -7989 -2460
rect -7969 2460 -2670 2600
rect -7969 -2460 -7749 2460
rect -2890 -2460 -2670 2460
rect -7969 -2600 -2670 -2460
rect -2650 2460 2649 2600
rect -2650 -2460 -2430 2460
rect 2429 -2460 2649 2460
rect -2650 -2600 2649 -2460
rect 2669 2460 7968 2600
rect 2669 -2460 2889 2460
rect 7748 -2460 7968 2460
rect 2669 -2600 7968 -2460
rect 7988 2460 13287 2600
rect 7988 -2460 8208 2460
rect 7988 -2600 13287 -2460
rect -13288 -2840 -7989 -2700
rect -8209 -7760 -7989 -2840
rect -13288 -7900 -7989 -7760
rect -7969 -2840 -2670 -2700
rect -7969 -7760 -7749 -2840
rect -2890 -7760 -2670 -2840
rect -7969 -7900 -2670 -7760
rect -2650 -2840 2649 -2700
rect -2650 -7760 -2430 -2840
rect 2429 -7760 2649 -2840
rect -2650 -7900 2649 -7760
rect 2669 -2840 7968 -2700
rect 2669 -7760 2889 -2840
rect 7748 -7760 7968 -2840
rect 2669 -7900 7968 -7760
rect 7988 -2840 13287 -2700
rect 7988 -7760 8208 -2840
rect 7988 -7900 13287 -7760
rect -13288 -8140 -7989 -8000
rect -8209 -13200 -7989 -8140
rect -7969 -8140 -2670 -8000
rect -7969 -13200 -7749 -8140
rect -2890 -13200 -2670 -8140
rect -2650 -8140 2649 -8000
rect -2650 -13200 -2430 -8140
rect 2429 -13200 2649 -8140
rect 2669 -8140 7968 -8000
rect 2669 -13200 2889 -8140
rect 7748 -13200 7968 -8140
rect 7988 -8140 13287 -8000
rect 7988 -13200 8208 -8140
<< metal3 >>
rect -13288 13172 -7989 13200
rect -13288 8028 -8073 13172
rect -8009 8028 -7989 13172
rect -13288 8000 -7989 8028
rect -7969 13172 -2670 13200
rect -7969 8028 -2754 13172
rect -2690 8028 -2670 13172
rect -7969 8000 -2670 8028
rect -2650 13172 2649 13200
rect -2650 8028 2565 13172
rect 2629 8028 2649 13172
rect -2650 8000 2649 8028
rect 2669 13172 7968 13200
rect 2669 8028 7884 13172
rect 7948 8028 7968 13172
rect 2669 8000 7968 8028
rect 7988 13172 13287 13200
rect 7988 8028 13203 13172
rect 13267 8028 13287 13172
rect 7988 8000 13287 8028
rect -13288 7872 -7989 7900
rect -13288 2728 -8073 7872
rect -8009 2728 -7989 7872
rect -13288 2700 -7989 2728
rect -7969 7872 -2670 7900
rect -7969 2728 -2754 7872
rect -2690 2728 -2670 7872
rect -7969 2700 -2670 2728
rect -2650 7872 2649 7900
rect -2650 2728 2565 7872
rect 2629 2728 2649 7872
rect -2650 2700 2649 2728
rect 2669 7872 7968 7900
rect 2669 2728 7884 7872
rect 7948 2728 7968 7872
rect 2669 2700 7968 2728
rect 7988 7872 13287 7900
rect 7988 2728 13203 7872
rect 13267 2728 13287 7872
rect 7988 2700 13287 2728
rect -13288 2572 -7989 2600
rect -13288 -2572 -8073 2572
rect -8009 -2572 -7989 2572
rect -13288 -2600 -7989 -2572
rect -7969 2572 -2670 2600
rect -7969 -2572 -2754 2572
rect -2690 -2572 -2670 2572
rect -7969 -2600 -2670 -2572
rect -2650 2572 2649 2600
rect -2650 -2572 2565 2572
rect 2629 -2572 2649 2572
rect -2650 -2600 2649 -2572
rect 2669 2572 7968 2600
rect 2669 -2572 7884 2572
rect 7948 -2572 7968 2572
rect 2669 -2600 7968 -2572
rect 7988 2572 13287 2600
rect 7988 -2572 13203 2572
rect 13267 -2572 13287 2572
rect 7988 -2600 13287 -2572
rect -13288 -2728 -7989 -2700
rect -13288 -7872 -8073 -2728
rect -8009 -7872 -7989 -2728
rect -13288 -7900 -7989 -7872
rect -7969 -2728 -2670 -2700
rect -7969 -7872 -2754 -2728
rect -2690 -7872 -2670 -2728
rect -7969 -7900 -2670 -7872
rect -2650 -2728 2649 -2700
rect -2650 -7872 2565 -2728
rect 2629 -7872 2649 -2728
rect -2650 -7900 2649 -7872
rect 2669 -2728 7968 -2700
rect 2669 -7872 7884 -2728
rect 7948 -7872 7968 -2728
rect 2669 -7900 7968 -7872
rect 7988 -2728 13287 -2700
rect 7988 -7872 13203 -2728
rect 13267 -7872 13287 -2728
rect 7988 -7900 13287 -7872
rect -13288 -8028 -7989 -8000
rect -13288 -13172 -8073 -8028
rect -8009 -13172 -7989 -8028
rect -13288 -13200 -7989 -13172
rect -7969 -8028 -2670 -8000
rect -7969 -13172 -2754 -8028
rect -2690 -13172 -2670 -8028
rect -7969 -13200 -2670 -13172
rect -2650 -8028 2649 -8000
rect -2650 -13172 2565 -8028
rect 2629 -13172 2649 -8028
rect -2650 -13200 2649 -13172
rect 2669 -8028 7968 -8000
rect 2669 -13172 7884 -8028
rect 7948 -13172 7968 -8028
rect 2669 -13200 7968 -13172
rect 7988 -8028 13287 -8000
rect 7988 -13172 13203 -8028
rect 13267 -13172 13287 -8028
rect 7988 -13200 13287 -13172
<< via3 >>
rect -8073 8028 -8009 13172
rect -2754 8028 -2690 13172
rect 2565 8028 2629 13172
rect 7884 8028 7948 13172
rect 13203 8028 13267 13172
rect -8073 2728 -8009 7872
rect -2754 2728 -2690 7872
rect 2565 2728 2629 7872
rect 7884 2728 7948 7872
rect 13203 2728 13267 7872
rect -8073 -2572 -8009 2572
rect -2754 -2572 -2690 2572
rect 2565 -2572 2629 2572
rect 7884 -2572 7948 2572
rect 13203 -2572 13267 2572
rect -8073 -7872 -8009 -2728
rect -2754 -7872 -2690 -2728
rect 2565 -7872 2629 -2728
rect 7884 -7872 7948 -2728
rect 13203 -7872 13267 -2728
rect -8073 -13172 -8009 -8028
rect -2754 -13172 -2690 -8028
rect 2565 -13172 2629 -8028
rect 7884 -13172 7948 -8028
rect 13203 -13172 13267 -8028
<< mimcap >>
rect -13188 13060 -8188 13100
rect -13188 8140 -13148 13060
rect -8228 8140 -8188 13060
rect -13188 8100 -8188 8140
rect -7869 13060 -2869 13100
rect -7869 8140 -7829 13060
rect -2909 8140 -2869 13060
rect -7869 8100 -2869 8140
rect -2550 13060 2450 13100
rect -2550 8140 -2510 13060
rect 2410 8140 2450 13060
rect -2550 8100 2450 8140
rect 2769 13060 7769 13100
rect 2769 8140 2809 13060
rect 7729 8140 7769 13060
rect 2769 8100 7769 8140
rect 8088 13060 13088 13100
rect 8088 8140 8128 13060
rect 13048 8140 13088 13060
rect 8088 8100 13088 8140
rect -13188 7760 -8188 7800
rect -13188 2840 -13148 7760
rect -8228 2840 -8188 7760
rect -13188 2800 -8188 2840
rect -7869 7760 -2869 7800
rect -7869 2840 -7829 7760
rect -2909 2840 -2869 7760
rect -7869 2800 -2869 2840
rect -2550 7760 2450 7800
rect -2550 2840 -2510 7760
rect 2410 2840 2450 7760
rect -2550 2800 2450 2840
rect 2769 7760 7769 7800
rect 2769 2840 2809 7760
rect 7729 2840 7769 7760
rect 2769 2800 7769 2840
rect 8088 7760 13088 7800
rect 8088 2840 8128 7760
rect 13048 2840 13088 7760
rect 8088 2800 13088 2840
rect -13188 2460 -8188 2500
rect -13188 -2460 -13148 2460
rect -8228 -2460 -8188 2460
rect -13188 -2500 -8188 -2460
rect -7869 2460 -2869 2500
rect -7869 -2460 -7829 2460
rect -2909 -2460 -2869 2460
rect -7869 -2500 -2869 -2460
rect -2550 2460 2450 2500
rect -2550 -2460 -2510 2460
rect 2410 -2460 2450 2460
rect -2550 -2500 2450 -2460
rect 2769 2460 7769 2500
rect 2769 -2460 2809 2460
rect 7729 -2460 7769 2460
rect 2769 -2500 7769 -2460
rect 8088 2460 13088 2500
rect 8088 -2460 8128 2460
rect 13048 -2460 13088 2460
rect 8088 -2500 13088 -2460
rect -13188 -2840 -8188 -2800
rect -13188 -7760 -13148 -2840
rect -8228 -7760 -8188 -2840
rect -13188 -7800 -8188 -7760
rect -7869 -2840 -2869 -2800
rect -7869 -7760 -7829 -2840
rect -2909 -7760 -2869 -2840
rect -7869 -7800 -2869 -7760
rect -2550 -2840 2450 -2800
rect -2550 -7760 -2510 -2840
rect 2410 -7760 2450 -2840
rect -2550 -7800 2450 -7760
rect 2769 -2840 7769 -2800
rect 2769 -7760 2809 -2840
rect 7729 -7760 7769 -2840
rect 2769 -7800 7769 -7760
rect 8088 -2840 13088 -2800
rect 8088 -7760 8128 -2840
rect 13048 -7760 13088 -2840
rect 8088 -7800 13088 -7760
rect -13188 -8140 -8188 -8100
rect -13188 -13060 -13148 -8140
rect -8228 -13060 -8188 -8140
rect -13188 -13100 -8188 -13060
rect -7869 -8140 -2869 -8100
rect -7869 -13060 -7829 -8140
rect -2909 -13060 -2869 -8140
rect -7869 -13100 -2869 -13060
rect -2550 -8140 2450 -8100
rect -2550 -13060 -2510 -8140
rect 2410 -13060 2450 -8140
rect -2550 -13100 2450 -13060
rect 2769 -8140 7769 -8100
rect 2769 -13060 2809 -8140
rect 7729 -13060 7769 -8140
rect 2769 -13100 7769 -13060
rect 8088 -8140 13088 -8100
rect 8088 -13060 8128 -8140
rect 13048 -13060 13088 -8140
rect 8088 -13100 13088 -13060
<< mimcapcontact >>
rect -13148 8140 -8228 13060
rect -7829 8140 -2909 13060
rect -2510 8140 2410 13060
rect 2809 8140 7729 13060
rect 8128 8140 13048 13060
rect -13148 2840 -8228 7760
rect -7829 2840 -2909 7760
rect -2510 2840 2410 7760
rect 2809 2840 7729 7760
rect 8128 2840 13048 7760
rect -13148 -2460 -8228 2460
rect -7829 -2460 -2909 2460
rect -2510 -2460 2410 2460
rect 2809 -2460 7729 2460
rect 8128 -2460 13048 2460
rect -13148 -7760 -8228 -2840
rect -7829 -7760 -2909 -2840
rect -2510 -7760 2410 -2840
rect 2809 -7760 7729 -2840
rect 8128 -7760 13048 -2840
rect -13148 -13060 -8228 -8140
rect -7829 -13060 -2909 -8140
rect -2510 -13060 2410 -8140
rect 2809 -13060 7729 -8140
rect 8128 -13060 13048 -8140
<< metal4 >>
rect -10740 13061 -10636 13250
rect -8120 13188 -8016 13250
rect -8120 13172 -7993 13188
rect -13149 13060 -8227 13061
rect -13149 8140 -13148 13060
rect -8228 8140 -8227 13060
rect -13149 8139 -8227 8140
rect -10740 7761 -10636 8139
rect -8120 8028 -8073 13172
rect -8009 8028 -7993 13172
rect -5421 13061 -5317 13250
rect -2801 13188 -2697 13250
rect -2801 13172 -2674 13188
rect -7830 13060 -2908 13061
rect -7830 8140 -7829 13060
rect -2909 8140 -2908 13060
rect -7830 8139 -2908 8140
rect -8120 8012 -7993 8028
rect -8120 7888 -8016 8012
rect -8120 7872 -7993 7888
rect -13149 7760 -8227 7761
rect -13149 2840 -13148 7760
rect -8228 2840 -8227 7760
rect -13149 2839 -8227 2840
rect -10740 2461 -10636 2839
rect -8120 2728 -8073 7872
rect -8009 2728 -7993 7872
rect -5421 7761 -5317 8139
rect -2801 8028 -2754 13172
rect -2690 8028 -2674 13172
rect -102 13061 2 13250
rect 2518 13188 2622 13250
rect 2518 13172 2645 13188
rect -2511 13060 2411 13061
rect -2511 8140 -2510 13060
rect 2410 8140 2411 13060
rect -2511 8139 2411 8140
rect -2801 8012 -2674 8028
rect -2801 7888 -2697 8012
rect -2801 7872 -2674 7888
rect -7830 7760 -2908 7761
rect -7830 2840 -7829 7760
rect -2909 2840 -2908 7760
rect -7830 2839 -2908 2840
rect -8120 2712 -7993 2728
rect -8120 2588 -8016 2712
rect -8120 2572 -7993 2588
rect -13149 2460 -8227 2461
rect -13149 -2460 -13148 2460
rect -8228 -2460 -8227 2460
rect -13149 -2461 -8227 -2460
rect -10740 -2839 -10636 -2461
rect -8120 -2572 -8073 2572
rect -8009 -2572 -7993 2572
rect -5421 2461 -5317 2839
rect -2801 2728 -2754 7872
rect -2690 2728 -2674 7872
rect -102 7761 2 8139
rect 2518 8028 2565 13172
rect 2629 8028 2645 13172
rect 5217 13061 5321 13250
rect 7837 13188 7941 13250
rect 7837 13172 7964 13188
rect 2808 13060 7730 13061
rect 2808 8140 2809 13060
rect 7729 8140 7730 13060
rect 2808 8139 7730 8140
rect 2518 8012 2645 8028
rect 2518 7888 2622 8012
rect 2518 7872 2645 7888
rect -2511 7760 2411 7761
rect -2511 2840 -2510 7760
rect 2410 2840 2411 7760
rect -2511 2839 2411 2840
rect -2801 2712 -2674 2728
rect -2801 2588 -2697 2712
rect -2801 2572 -2674 2588
rect -7830 2460 -2908 2461
rect -7830 -2460 -7829 2460
rect -2909 -2460 -2908 2460
rect -7830 -2461 -2908 -2460
rect -8120 -2588 -7993 -2572
rect -8120 -2712 -8016 -2588
rect -8120 -2728 -7993 -2712
rect -13149 -2840 -8227 -2839
rect -13149 -7760 -13148 -2840
rect -8228 -7760 -8227 -2840
rect -13149 -7761 -8227 -7760
rect -10740 -8139 -10636 -7761
rect -8120 -7872 -8073 -2728
rect -8009 -7872 -7993 -2728
rect -5421 -2839 -5317 -2461
rect -2801 -2572 -2754 2572
rect -2690 -2572 -2674 2572
rect -102 2461 2 2839
rect 2518 2728 2565 7872
rect 2629 2728 2645 7872
rect 5217 7761 5321 8139
rect 7837 8028 7884 13172
rect 7948 8028 7964 13172
rect 10536 13061 10640 13250
rect 13156 13188 13260 13250
rect 13156 13172 13283 13188
rect 8127 13060 13049 13061
rect 8127 8140 8128 13060
rect 13048 8140 13049 13060
rect 8127 8139 13049 8140
rect 7837 8012 7964 8028
rect 7837 7888 7941 8012
rect 7837 7872 7964 7888
rect 2808 7760 7730 7761
rect 2808 2840 2809 7760
rect 7729 2840 7730 7760
rect 2808 2839 7730 2840
rect 2518 2712 2645 2728
rect 2518 2588 2622 2712
rect 2518 2572 2645 2588
rect -2511 2460 2411 2461
rect -2511 -2460 -2510 2460
rect 2410 -2460 2411 2460
rect -2511 -2461 2411 -2460
rect -2801 -2588 -2674 -2572
rect -2801 -2712 -2697 -2588
rect -2801 -2728 -2674 -2712
rect -7830 -2840 -2908 -2839
rect -7830 -7760 -7829 -2840
rect -2909 -7760 -2908 -2840
rect -7830 -7761 -2908 -7760
rect -8120 -7888 -7993 -7872
rect -8120 -8012 -8016 -7888
rect -8120 -8028 -7993 -8012
rect -13149 -8140 -8227 -8139
rect -13149 -13060 -13148 -8140
rect -8228 -13060 -8227 -8140
rect -13149 -13061 -8227 -13060
rect -10740 -13250 -10636 -13061
rect -8120 -13172 -8073 -8028
rect -8009 -13172 -7993 -8028
rect -5421 -8139 -5317 -7761
rect -2801 -7872 -2754 -2728
rect -2690 -7872 -2674 -2728
rect -102 -2839 2 -2461
rect 2518 -2572 2565 2572
rect 2629 -2572 2645 2572
rect 5217 2461 5321 2839
rect 7837 2728 7884 7872
rect 7948 2728 7964 7872
rect 10536 7761 10640 8139
rect 13156 8028 13203 13172
rect 13267 8028 13283 13172
rect 13156 8012 13283 8028
rect 13156 7888 13260 8012
rect 13156 7872 13283 7888
rect 8127 7760 13049 7761
rect 8127 2840 8128 7760
rect 13048 2840 13049 7760
rect 8127 2839 13049 2840
rect 7837 2712 7964 2728
rect 7837 2588 7941 2712
rect 7837 2572 7964 2588
rect 2808 2460 7730 2461
rect 2808 -2460 2809 2460
rect 7729 -2460 7730 2460
rect 2808 -2461 7730 -2460
rect 2518 -2588 2645 -2572
rect 2518 -2712 2622 -2588
rect 2518 -2728 2645 -2712
rect -2511 -2840 2411 -2839
rect -2511 -7760 -2510 -2840
rect 2410 -7760 2411 -2840
rect -2511 -7761 2411 -7760
rect -2801 -7888 -2674 -7872
rect -2801 -8012 -2697 -7888
rect -2801 -8028 -2674 -8012
rect -7830 -8140 -2908 -8139
rect -7830 -13060 -7829 -8140
rect -2909 -13060 -2908 -8140
rect -7830 -13061 -2908 -13060
rect -8120 -13188 -7993 -13172
rect -8120 -13250 -8016 -13188
rect -5421 -13250 -5317 -13061
rect -2801 -13172 -2754 -8028
rect -2690 -13172 -2674 -8028
rect -102 -8139 2 -7761
rect 2518 -7872 2565 -2728
rect 2629 -7872 2645 -2728
rect 5217 -2839 5321 -2461
rect 7837 -2572 7884 2572
rect 7948 -2572 7964 2572
rect 10536 2461 10640 2839
rect 13156 2728 13203 7872
rect 13267 2728 13283 7872
rect 13156 2712 13283 2728
rect 13156 2588 13260 2712
rect 13156 2572 13283 2588
rect 8127 2460 13049 2461
rect 8127 -2460 8128 2460
rect 13048 -2460 13049 2460
rect 8127 -2461 13049 -2460
rect 7837 -2588 7964 -2572
rect 7837 -2712 7941 -2588
rect 7837 -2728 7964 -2712
rect 2808 -2840 7730 -2839
rect 2808 -7760 2809 -2840
rect 7729 -7760 7730 -2840
rect 2808 -7761 7730 -7760
rect 2518 -7888 2645 -7872
rect 2518 -8012 2622 -7888
rect 2518 -8028 2645 -8012
rect -2511 -8140 2411 -8139
rect -2511 -13060 -2510 -8140
rect 2410 -13060 2411 -8140
rect -2511 -13061 2411 -13060
rect -2801 -13188 -2674 -13172
rect -2801 -13250 -2697 -13188
rect -102 -13250 2 -13061
rect 2518 -13172 2565 -8028
rect 2629 -13172 2645 -8028
rect 5217 -8139 5321 -7761
rect 7837 -7872 7884 -2728
rect 7948 -7872 7964 -2728
rect 10536 -2839 10640 -2461
rect 13156 -2572 13203 2572
rect 13267 -2572 13283 2572
rect 13156 -2588 13283 -2572
rect 13156 -2712 13260 -2588
rect 13156 -2728 13283 -2712
rect 8127 -2840 13049 -2839
rect 8127 -7760 8128 -2840
rect 13048 -7760 13049 -2840
rect 8127 -7761 13049 -7760
rect 7837 -7888 7964 -7872
rect 7837 -8012 7941 -7888
rect 7837 -8028 7964 -8012
rect 2808 -8140 7730 -8139
rect 2808 -13060 2809 -8140
rect 7729 -13060 7730 -8140
rect 2808 -13061 7730 -13060
rect 2518 -13188 2645 -13172
rect 2518 -13250 2622 -13188
rect 5217 -13250 5321 -13061
rect 7837 -13172 7884 -8028
rect 7948 -13172 7964 -8028
rect 10536 -8139 10640 -7761
rect 13156 -7872 13203 -2728
rect 13267 -7872 13283 -2728
rect 13156 -7888 13283 -7872
rect 13156 -8012 13260 -7888
rect 13156 -8028 13283 -8012
rect 8127 -8140 13049 -8139
rect 8127 -13060 8128 -8140
rect 13048 -13060 13049 -8140
rect 8127 -13061 13049 -13060
rect 7837 -13188 7964 -13172
rect 7837 -13250 7941 -13188
rect 10536 -13250 10640 -13061
rect 13156 -13172 13203 -8028
rect 13267 -13172 13283 -8028
rect 13156 -13188 13283 -13172
rect 13156 -13250 13260 -13188
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 7988 8000 13188 13200
string parameters w 25 l 25 val 1.269k carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
