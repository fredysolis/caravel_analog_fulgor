magic
tech sky130A
magscale 1 2
timestamp 1623451718
<< pwell >>
rect -263 -255 263 255
<< nmos >>
rect -63 -45 -33 45
rect 33 -45 63 45
<< ndiff >>
rect -125 33 -63 45
rect -125 -33 -113 33
rect -79 -33 -63 33
rect -125 -45 -63 -33
rect -33 33 33 45
rect -33 -33 -17 33
rect 17 -33 33 33
rect -33 -45 33 -33
rect 63 33 125 45
rect 63 -33 79 33
rect 113 -33 125 33
rect 63 -45 125 -33
<< ndiffc >>
rect -113 -33 -79 33
rect -17 -33 17 33
rect 79 -33 113 33
<< psubdiff >>
rect -193 -219 -131 -185
rect 131 -219 193 -185
<< psubdiffcont >>
rect -131 -219 131 -185
<< poly >>
rect -129 71 -33 137
rect -63 45 -33 71
rect 33 67 99 133
rect 33 45 63 67
rect -63 -71 -33 -45
rect 33 -71 63 -45
<< locali >>
rect -113 33 -79 49
rect -113 -49 -79 -33
rect -17 33 17 49
rect -17 -49 17 -33
rect 79 33 113 49
rect 79 -49 113 -33
rect -193 -219 -131 -185
rect 131 -219 193 -185
<< viali >>
rect -113 -33 -79 33
rect -17 -33 17 33
rect 79 -33 113 33
<< metal1 >>
rect -119 33 -73 45
rect -119 -33 -113 33
rect -79 -33 -73 33
rect -119 -45 -73 -33
rect -23 33 23 45
rect -23 -33 -17 33
rect 17 -33 23 33
rect -23 -45 23 -33
rect 73 33 119 45
rect 73 -33 79 33
rect 113 -33 119 33
rect 73 -45 119 -33
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -210 -202 210 202
string parameters w 0.45 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
