magic
tech sky130A
magscale 1 2
timestamp 1623958459
<< pwell >>
rect -551 188 551 310
rect -551 122 -302 188
rect -298 122 -178 188
rect -176 122 274 188
rect 277 122 551 188
rect -551 -310 551 122
<< nmoslvt >>
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
<< ndiff >>
rect -413 88 -351 100
rect -413 -88 -401 88
rect -367 -88 -351 88
rect -413 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 413 100
rect 351 -88 367 88
rect 401 -88 413 88
rect 351 -100 413 -88
<< ndiffc >>
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
<< psubdiff >>
rect -515 240 -419 274
rect 419 240 515 274
rect -515 178 -481 240
rect 481 178 515 240
rect -515 -240 -481 -178
rect 481 -240 515 -178
rect -515 -274 -419 -240
rect 419 -274 515 -240
<< psubdiffcont >>
rect -419 240 419 274
rect -515 -178 -481 178
rect 481 -178 515 178
rect -419 -274 419 -240
<< poly >>
rect -368 172 369 188
rect -368 138 -352 172
rect -318 138 -257 172
rect -223 138 -160 172
rect -126 138 -65 172
rect -31 138 32 172
rect 66 138 127 172
rect 161 138 224 172
rect 258 138 319 172
rect 353 138 369 172
rect -368 122 369 138
rect -351 100 -321 122
rect -255 100 -225 122
rect -159 100 -129 122
rect -63 100 -33 122
rect 33 100 63 122
rect 129 100 159 122
rect 225 100 255 122
rect 321 100 351 122
rect -351 -126 -321 -100
rect -255 -126 -225 -100
rect -159 -126 -129 -100
rect -63 -126 -33 -100
rect 33 -126 63 -100
rect 129 -126 159 -100
rect 225 -126 255 -100
rect 321 -126 351 -100
<< polycont >>
rect -352 138 -318 172
rect -257 138 -223 172
rect -160 138 -126 172
rect -65 138 -31 172
rect 32 138 66 172
rect 127 138 161 172
rect 224 138 258 172
rect 319 138 353 172
<< locali >>
rect -515 240 -419 274
rect 419 240 515 274
rect -515 178 -481 240
rect 481 178 515 240
rect -368 138 -352 172
rect 353 138 369 172
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect -515 -240 -481 -178
rect 481 -240 515 -178
rect -515 -274 -419 -240
rect 419 -274 515 -240
<< viali >>
rect -352 138 -318 172
rect -318 138 -257 172
rect -257 138 -223 172
rect -223 138 -160 172
rect -160 138 -126 172
rect -126 138 -65 172
rect -65 138 -31 172
rect -31 138 32 172
rect 32 138 66 172
rect 66 138 127 172
rect 127 138 161 172
rect 161 138 224 172
rect 224 138 258 172
rect 258 138 319 172
rect 319 138 353 172
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
<< metal1 >>
rect -364 172 365 178
rect -364 138 -352 172
rect 353 138 365 172
rect -364 132 365 138
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -498 -257 498 257
string parameters w 1 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
