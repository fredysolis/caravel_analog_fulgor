magic
tech sky130A
magscale 1 2
timestamp 1624020979
<< nwell >>
rect -263 -319 263 319
<< pmos >>
rect -63 -100 -33 100
rect 33 -100 63 100
<< pdiff >>
rect -125 88 -63 100
rect -125 -88 -113 88
rect -79 -88 -63 88
rect -125 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 125 100
rect 63 -88 79 88
rect 113 -88 125 88
rect 63 -100 125 -88
<< pdiffc >>
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
<< nsubdiff >>
rect -227 249 -131 283
rect 131 249 227 283
rect -227 187 -193 249
rect 193 187 227 249
rect -227 -249 -193 -187
rect 193 -249 227 -187
rect -227 -283 -131 -249
rect 131 -283 227 -249
<< nsubdiffcont >>
rect -131 249 131 283
rect -227 -187 -193 187
rect 193 -187 227 187
rect -131 -283 131 -249
<< poly >>
rect -63 100 -33 126
rect 33 100 63 126
rect -63 -131 -33 -100
rect 33 -131 63 -100
rect -81 -147 81 -131
rect -81 -181 -65 -147
rect -31 -181 31 -147
rect 65 -181 81 -147
rect -81 -197 81 -181
<< polycont >>
rect -65 -181 -31 -147
rect 31 -181 65 -147
<< locali >>
rect -227 249 -131 283
rect 131 249 227 283
rect -227 187 -193 249
rect 193 187 227 249
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect -81 -181 -65 -147
rect -31 -181 31 -147
rect 65 -181 81 -147
rect -227 -249 -193 -187
rect 193 -249 227 -187
rect -227 -283 -131 -249
rect 131 -283 227 -249
<< viali >>
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect -65 -181 -31 -147
rect 31 -181 65 -147
<< metal1 >>
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect -77 -147 77 -141
rect -77 -181 -65 -147
rect -31 -181 31 -147
rect 65 -181 77 -147
rect -77 -187 77 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -210 -266 210 266
string parameters w 1 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
