**.subckt mux2to4 in_a in_b selec_0_neg selec_0 out_b_0 out_b_1 out_a_0 out_a_1 vdd vss
*.iopin in_a
*.iopin in_b
*.ipin selec_0_neg
*.ipin selec_0
*.iopin out_b_0
*.iopin out_b_1
*.iopin out_a_0
*.iopin out_a_1
*.iopin vdd
*.iopin vss
x4 selec_0 out_a_1 in_a selec_0_neg vss vdd trans_gate_mux2to8
x5 selec_0_neg out_a_0 in_a selec_0 vss vdd trans_gate_mux2to8
x8 selec_0 out_b_1 in_b selec_0_neg vss vdd trans_gate_mux2to8
x9 selec_0_neg out_b_0 in_b selec_0 vss vdd trans_gate_mux2to8
**.ends

* expanding   symbol:  trans_gate_mux2to8.sym # of pins=6
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/trans_gate_mux2to8.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/trans_gate_mux2to8.sch
.subckt trans_gate_mux2to8  en_pos out in en_neg vss vdd
*.iopin en_neg
*.ipin in
*.opin out
*.iopin en_pos
*.iopin vdd
*.iopin vss
XM2 out en_neg in vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM1 out en_pos in vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
.ends

** flattened .save nodes
.end
