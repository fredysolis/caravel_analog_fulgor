magic
tech sky130A
magscale 1 2
timestamp 1623976832
<< nwell >>
rect -807 -384 807 384
<< pmoslvt >>
rect -611 -236 -541 164
rect -483 -236 -413 164
rect -355 -236 -285 164
rect -227 -236 -157 164
rect -99 -236 -29 164
rect 29 -236 99 164
rect 157 -236 227 164
rect 285 -236 355 164
rect 413 -236 483 164
rect 541 -236 611 164
<< pdiff >>
rect -669 152 -611 164
rect -669 -224 -657 152
rect -623 -224 -611 152
rect -669 -236 -611 -224
rect -541 152 -483 164
rect -541 -224 -529 152
rect -495 -224 -483 152
rect -541 -236 -483 -224
rect -413 152 -355 164
rect -413 -224 -401 152
rect -367 -224 -355 152
rect -413 -236 -355 -224
rect -285 152 -227 164
rect -285 -224 -273 152
rect -239 -224 -227 152
rect -285 -236 -227 -224
rect -157 152 -99 164
rect -157 -224 -145 152
rect -111 -224 -99 152
rect -157 -236 -99 -224
rect -29 152 29 164
rect -29 -224 -17 152
rect 17 -224 29 152
rect -29 -236 29 -224
rect 99 152 157 164
rect 99 -224 111 152
rect 145 -224 157 152
rect 99 -236 157 -224
rect 227 152 285 164
rect 227 -224 239 152
rect 273 -224 285 152
rect 227 -236 285 -224
rect 355 152 413 164
rect 355 -224 367 152
rect 401 -224 413 152
rect 355 -236 413 -224
rect 483 152 541 164
rect 483 -224 495 152
rect 529 -224 541 152
rect 483 -236 541 -224
rect 611 152 669 164
rect 611 -224 623 152
rect 657 -224 669 152
rect 611 -236 669 -224
<< pdiffc >>
rect -657 -224 -623 152
rect -529 -224 -495 152
rect -401 -224 -367 152
rect -273 -224 -239 152
rect -145 -224 -111 152
rect -17 -224 17 152
rect 111 -224 145 152
rect 239 -224 273 152
rect 367 -224 401 152
rect 495 -224 529 152
rect 623 -224 657 152
<< nsubdiff >>
rect -771 314 -675 348
rect 675 314 771 348
rect -771 251 -737 314
rect 737 251 771 314
rect -771 -314 -737 -251
rect 737 -314 771 -251
rect -771 -348 -675 -314
rect 675 -348 771 -314
<< nsubdiffcont >>
rect -675 314 675 348
rect -771 -251 -737 251
rect 737 -251 771 251
rect -675 -348 675 -314
<< poly >>
rect -611 245 611 261
rect -611 211 -595 245
rect -557 211 -467 245
rect -429 211 -339 245
rect -301 211 -211 245
rect -173 211 -83 245
rect -45 211 45 245
rect 83 211 173 245
rect 211 211 301 245
rect 339 211 429 245
rect 467 211 557 245
rect 595 211 611 245
rect -611 201 611 211
rect -611 164 -541 201
rect -483 164 -413 201
rect -355 164 -285 201
rect -227 164 -157 201
rect -99 164 -29 201
rect 29 164 99 201
rect 157 164 227 201
rect 285 164 355 201
rect 413 164 483 201
rect 541 164 611 201
rect -611 -262 -541 -236
rect -483 -262 -413 -236
rect -355 -262 -285 -236
rect -227 -262 -157 -236
rect -99 -262 -29 -236
rect 29 -262 99 -236
rect 157 -262 227 -236
rect 285 -262 355 -236
rect 413 -262 483 -236
rect 541 -262 611 -236
<< polycont >>
rect -595 211 -557 245
rect -467 211 -429 245
rect -339 211 -301 245
rect -211 211 -173 245
rect -83 211 -45 245
rect 45 211 83 245
rect 173 211 211 245
rect 301 211 339 245
rect 429 211 467 245
rect 557 211 595 245
<< locali >>
rect -771 314 -675 348
rect 675 314 771 348
rect -771 251 -737 314
rect 737 251 771 314
rect -611 211 -595 245
rect 595 211 611 245
rect -657 152 -623 168
rect -657 -240 -623 -224
rect -529 152 -495 168
rect -529 -240 -495 -224
rect -401 152 -367 168
rect -401 -240 -367 -224
rect -273 152 -239 168
rect -273 -240 -239 -224
rect -145 152 -111 168
rect -145 -240 -111 -224
rect -17 152 17 168
rect -17 -240 17 -224
rect 111 152 145 168
rect 111 -240 145 -224
rect 239 152 273 168
rect 239 -240 273 -224
rect 367 152 401 168
rect 367 -240 401 -224
rect 495 152 529 168
rect 495 -240 529 -224
rect 623 152 657 168
rect 623 -240 657 -224
rect -771 -314 -737 -251
rect 737 -314 771 -251
rect -771 -348 -675 -314
rect 675 -348 771 -314
<< viali >>
rect -595 211 -557 245
rect -557 211 -467 245
rect -467 211 -429 245
rect -429 211 -339 245
rect -339 211 -301 245
rect -301 211 -211 245
rect -211 211 -173 245
rect -173 211 -83 245
rect -83 211 -45 245
rect -45 211 45 245
rect 45 211 83 245
rect 83 211 173 245
rect 173 211 211 245
rect 211 211 301 245
rect 301 211 339 245
rect 339 211 429 245
rect 429 211 467 245
rect 467 211 557 245
rect 557 211 595 245
rect -657 -224 -623 152
rect -529 -224 -495 152
rect -401 -224 -367 152
rect -273 -224 -239 152
rect -145 -224 -111 152
rect -17 -224 17 152
rect 111 -224 145 152
rect 239 -224 273 152
rect 367 -224 401 152
rect 495 -224 529 152
rect 623 -224 657 152
<< metal1 >>
rect -607 245 607 251
rect -607 211 -595 245
rect 595 211 607 245
rect -607 205 607 211
rect -663 152 -617 164
rect -663 -224 -657 152
rect -623 -224 -617 152
rect -663 -236 -617 -224
rect -535 152 -489 164
rect -535 -224 -529 152
rect -495 -224 -489 152
rect -535 -236 -489 -224
rect -407 152 -361 164
rect -407 -224 -401 152
rect -367 -224 -361 152
rect -407 -236 -361 -224
rect -279 152 -233 164
rect -279 -224 -273 152
rect -239 -224 -233 152
rect -279 -236 -233 -224
rect -151 152 -105 164
rect -151 -224 -145 152
rect -111 -224 -105 152
rect -151 -236 -105 -224
rect -23 152 23 164
rect -23 -224 -17 152
rect 17 -224 23 152
rect -23 -236 23 -224
rect 105 152 151 164
rect 105 -224 111 152
rect 145 -224 151 152
rect 105 -236 151 -224
rect 233 152 279 164
rect 233 -224 239 152
rect 273 -224 279 152
rect 233 -236 279 -224
rect 361 152 407 164
rect 361 -224 367 152
rect 401 -224 407 152
rect 361 -236 407 -224
rect 489 152 535 164
rect 489 -224 495 152
rect 529 -224 535 152
rect 489 -236 535 -224
rect 617 152 663 164
rect 617 -224 623 152
rect 657 -224 663 152
rect 617 -236 663 -224
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -754 -331 754 331
string parameters w 2 l 0.35 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
