magic
tech sky130A
magscale 1 2
timestamp 1624395098
<< nwell >>
rect -556 2925 0 3068
rect -556 2664 57 2925
rect -111 2561 57 2664
rect -40 2555 57 2561
rect -30 2544 57 2555
rect 1803 2292 7702 3068
rect 9171 2292 9793 3068
rect 12155 2292 12777 3068
rect 13336 2664 13892 3068
rect -556 0 0 776
rect 1803 0 2425 776
rect 2984 0 3540 404
rect 5343 0 11242 776
rect 12155 0 12777 776
rect 13336 0 13892 776
<< pwell >>
rect -556 2241 -150 2292
rect -40 2241 0 2292
rect -556 776 0 2241
rect 5965 776 7368 2292
rect 13336 776 13892 2292
<< viali >>
rect -134 2343 -55 2507
rect 13765 2324 13836 2537
rect -312 2204 -237 2294
rect 6771 2238 7063 2299
rect 7175 2196 7309 2283
rect 13405 2206 13518 2260
rect 13581 2230 13645 2316
rect -523 2043 -356 2093
rect 6736 2050 6825 2183
rect 2989 974 3189 1025
rect 3228 773 3304 866
rect 3406 536 3486 738
<< metal1 >>
rect -556 2904 13892 3038
rect -357 2643 -199 2904
rect 6819 2643 7074 2904
rect 13535 2643 13693 2904
rect 13759 2537 13842 2549
rect -144 2330 -134 2521
rect -55 2330 -45 2521
rect -333 2199 -323 2317
rect -223 2199 -213 2317
rect 6263 2308 7075 2367
rect 6759 2299 7075 2308
rect 6759 2238 6771 2299
rect 7063 2238 7075 2299
rect 6759 2232 7075 2238
rect -318 2192 -231 2199
rect 7163 2196 7175 2336
rect 7309 2196 7321 2336
rect 13395 2266 13405 2298
rect 13393 2206 13405 2266
rect 13518 2266 13528 2298
rect 13518 2206 13530 2266
rect 13569 2230 13579 2334
rect 13645 2230 13655 2334
rect 13759 2324 13765 2537
rect 13836 2324 13842 2537
rect 13759 2312 13842 2324
rect 13575 2218 13651 2230
rect 13393 2200 13530 2206
rect -535 2093 -516 2152
rect -385 2093 -344 2152
rect 1987 2120 1997 2184
rect 2237 2120 2247 2184
rect 5527 2120 5537 2184
rect 5777 2120 5787 2184
rect 6730 2183 6831 2195
rect 7163 2190 7321 2196
rect -535 2043 -523 2093
rect -356 2043 -344 2093
rect 6701 2050 6711 2183
rect 6849 2050 6859 2183
rect 9355 2120 9365 2184
rect 9605 2120 9615 2184
rect 12339 2120 12349 2184
rect 12589 2120 12599 2184
rect -535 2037 -516 2043
rect -385 2037 -344 2043
rect 6730 2038 6831 2050
rect -357 1698 -199 1943
rect 6819 1698 7073 1944
rect 13535 1698 13693 1943
rect -556 1416 36 1698
rect -556 1370 0 1416
rect 2984 1370 3540 1698
rect 6524 1370 7371 1698
rect 13317 1370 13892 1698
rect 3183 1125 3341 1370
rect 2964 1025 3201 1031
rect 2964 974 2989 1025
rect 3189 974 3201 1025
rect 2964 968 3201 974
rect 1981 884 1991 948
rect 2231 884 2241 948
rect 2964 760 3023 968
rect 5521 884 5531 948
rect 5771 884 5781 948
rect 9349 884 9359 948
rect 9599 884 9609 948
rect 12333 884 12343 948
rect 12583 884 12593 948
rect 3222 872 3310 878
rect 3218 771 3228 872
rect 3304 771 3314 872
rect 3222 761 3310 771
rect 2652 701 3023 760
rect 3400 738 3492 750
rect 3396 536 3406 738
rect 3486 536 3496 738
rect 3400 524 3492 536
rect 3183 164 3341 425
rect -556 30 13892 164
<< via1 >>
rect -134 2507 -55 2521
rect -134 2343 -55 2507
rect -134 2330 -55 2343
rect -323 2294 -223 2317
rect -323 2204 -312 2294
rect -312 2204 -237 2294
rect -237 2204 -223 2294
rect -323 2199 -223 2204
rect 7175 2283 7309 2336
rect 7175 2196 7309 2283
rect 13405 2260 13518 2298
rect 13405 2206 13518 2260
rect 13579 2316 13645 2334
rect 13579 2230 13581 2316
rect 13581 2230 13645 2316
rect -516 2093 -385 2152
rect 1997 2120 2237 2184
rect 5537 2120 5777 2184
rect -516 2043 -385 2093
rect 6711 2050 6736 2183
rect 6736 2050 6825 2183
rect 6825 2050 6849 2183
rect 9365 2120 9605 2184
rect 12349 2120 12589 2184
rect -516 2037 -385 2043
rect 1991 884 2231 948
rect 5531 884 5771 948
rect 9359 884 9599 948
rect 12343 884 12583 948
rect 3228 866 3304 872
rect 3228 773 3304 866
rect 3228 771 3304 773
rect 3406 536 3486 738
<< metal2 >>
rect -516 2737 7309 2869
rect -516 2152 -384 2737
rect 7175 2700 7309 2737
rect -326 2568 6364 2700
rect -326 2317 -221 2568
rect -326 2199 -323 2317
rect -223 2199 -221 2317
rect -134 2521 -55 2531
rect -134 2254 227 2330
rect 6232 2287 6364 2568
rect 7175 2685 10684 2700
rect 7175 2573 10572 2685
rect 7175 2568 10684 2573
rect 7175 2336 7309 2568
rect 10572 2563 10684 2568
rect 13089 2464 13529 2540
rect -326 2197 -221 2199
rect -323 2189 -223 2197
rect 10137 2259 10572 2325
rect 13395 2298 13529 2464
rect 13395 2206 13405 2298
rect 13518 2206 13529 2298
rect 13395 2196 13529 2206
rect 13569 2230 13579 2334
rect 13645 2230 13655 2334
rect -385 2037 -384 2152
rect 1997 2184 2237 2194
rect 1997 2110 2237 2120
rect 5537 2184 5777 2194
rect 5537 2110 5777 2120
rect 6711 2183 6849 2193
rect 7175 2186 7309 2196
rect -516 2015 -384 2037
rect 9365 2184 9605 2194
rect 9365 2110 9605 2120
rect 12349 2184 12589 2194
rect 12349 2110 12589 2120
rect 6095 1601 6151 1611
rect 3237 1518 6095 1594
rect 1991 948 2231 958
rect 1991 874 2231 884
rect 3237 882 3313 1518
rect 6095 1469 6151 1479
rect 6711 1599 6849 2050
rect 6711 1591 7683 1599
rect 6711 1469 7617 1591
rect 7673 1469 7683 1591
rect 10133 1590 10189 1600
rect 10131 1498 10133 1570
rect 6711 1461 7683 1469
rect 10601 1590 10657 1600
rect 10189 1498 10601 1570
rect 10133 1468 10189 1478
rect 10657 1550 11273 1570
rect 13569 1564 13655 2230
rect 11484 1550 13655 1564
rect 10657 1478 13655 1550
rect 10601 1468 10657 1478
rect 3228 872 3313 882
rect 5531 948 5771 958
rect 5531 874 5771 884
rect 9359 948 9599 958
rect 9359 874 9599 884
rect 12343 948 12583 958
rect 12343 874 12583 884
rect 3304 776 3313 872
rect 3228 761 3304 771
rect 3406 738 3767 814
rect 10131 743 10578 809
rect 3406 526 3486 536
rect 3406 525 3482 526
<< via2 >>
rect 10572 2573 10684 2685
rect 1997 2120 2237 2184
rect 5537 2120 5777 2184
rect 9365 2120 9605 2184
rect 12349 2120 12589 2184
rect 1991 884 2231 948
rect 6095 1479 6151 1601
rect 7617 1469 7673 1591
rect 10133 1478 10189 1590
rect 10601 1478 10657 1590
rect 5531 884 5771 948
rect 9359 884 9599 948
rect 12343 884 12583 948
<< metal3 >>
rect 10562 2685 10694 2690
rect 10562 2573 10572 2685
rect 10684 2573 10694 2685
rect 10562 2568 10694 2573
rect 1987 2184 2247 2189
rect 1987 2120 1997 2184
rect 2237 2120 2247 2184
rect 1987 2115 2247 2120
rect 5527 2184 5787 2189
rect 5527 2120 5537 2184
rect 5777 2120 5787 2184
rect 5527 2115 5787 2120
rect 9355 2184 9615 2189
rect 9355 2120 9365 2184
rect 9605 2120 9615 2184
rect 9355 2115 9615 2120
rect 6085 1601 6161 1606
rect 6085 1479 6095 1601
rect 6151 1479 6161 1601
rect 6085 1474 6161 1479
rect 7607 1591 7683 1596
rect 10599 1595 10659 2568
rect 12339 2184 12599 2189
rect 12339 2120 12349 2184
rect 12589 2120 12599 2184
rect 12339 2115 12599 2120
rect 7607 1469 7617 1591
rect 7673 1469 7683 1591
rect 10123 1590 10199 1595
rect 10123 1478 10133 1590
rect 10189 1478 10199 1590
rect 10123 1473 10199 1478
rect 10591 1590 10667 1595
rect 10591 1478 10601 1590
rect 10657 1478 10667 1590
rect 10591 1473 10667 1478
rect 7607 1464 7683 1469
rect 1981 948 2241 953
rect 1981 884 1991 948
rect 2231 884 2241 948
rect 1981 879 2241 884
rect 5521 948 5781 953
rect 5521 884 5531 948
rect 5771 884 5781 948
rect 5521 879 5781 884
rect 9349 948 9609 953
rect 9349 884 9359 948
rect 9599 884 9609 948
rect 9349 879 9609 884
rect 10599 804 10659 1473
rect 12333 948 12593 953
rect 12333 884 12343 948
rect 12583 884 12593 948
rect 12333 879 12593 884
<< via3 >>
rect 1997 2120 2237 2184
rect 5537 2120 5777 2184
rect 9365 2120 9605 2184
rect 12349 2120 12589 2184
rect 1991 884 2231 948
rect 5531 884 5771 948
rect 9359 884 9599 948
rect 12343 884 12583 948
<< metal4 >>
rect 1996 2184 12590 2185
rect 1996 2120 1997 2184
rect 2237 2120 5537 2184
rect 5777 2120 9365 2184
rect 9605 2120 12349 2184
rect 12589 2120 12590 2184
rect 1996 2119 12590 2120
rect 1990 948 12584 949
rect 1990 884 1991 948
rect 2231 884 5531 948
rect 5771 884 9359 948
rect 9599 884 12343 948
rect 12583 884 12584 948
rect 1990 883 12584 884
use DFlipFlop  DFlipFlop_3
timestamp 1624049879
transform 1 0 11596 0 -1 3068
box -1244 0 1740 3068
use DFlipFlop  DFlipFlop_1
timestamp 1624049879
transform 1 0 4784 0 1 0
box -1244 0 1740 3068
use DFlipFlop  DFlipFlop_2
timestamp 1624049879
transform 1 0 8612 0 1 0
box -1244 0 1740 3068
use DFlipFlop  DFlipFlop_0
timestamp 1624049879
transform 1 0 1244 0 1 0
box -1244 0 1740 3068
use sky130_fd_sc_hs__or2_1  sky130_fd_sc_hs__or2_1_0
timestamp 1624049879
transform 1 0 13374 0 1 1960
box -38 -49 518 715
use sky130_fd_sc_hs__and2_1  sky130_fd_sc_hs__and2_1_0
timestamp 1624049879
transform 1 0 -518 0 1 1960
box -38 -49 518 715
use sky130_fd_sc_hs__xor2_1  sky130_fd_sc_hs__xor2_1_0
timestamp 1624049879
transform -1 0 7330 0 1 1960
box -38 -49 806 715
use sky130_fd_sc_hs__and2_1  sky130_fd_sc_hs__and2_1_1
timestamp 1624049879
transform 1 0 3022 0 -1 1108
box -38 -49 518 715
<< labels >>
rlabel metal2 7175 2568 10572 2700 1 Q1
rlabel metal1 6263 2308 7075 2367 1 Q0
rlabel metal1 -556 1370 0 1698 1 vss
rlabel metal1 2652 701 3023 760 1 nQ2
rlabel metal4 5771 883 9359 949 1 CLK
rlabel metal4 5777 2119 9365 2185 1 nCLK
rlabel metal1 -556 2904 13892 3038 1 vdd
rlabel viali 13765 2324 13836 2537 1 CLK_5
rlabel metal2 3237 1518 6095 1594 1 nQ0
rlabel metal2 13089 2464 13529 2540 1 Q1_shift
<< end >>
