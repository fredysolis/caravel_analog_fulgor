magic
tech sky130A
magscale 1 2
timestamp 1624885207
<< nwell >>
rect 2984 1980 4570 3060
rect 10382 2725 10536 3068
rect 10538 3058 10785 3068
rect 10538 2297 11706 3058
rect 10538 1971 11703 2297
rect 2984 1080 4332 1086
rect 2984 0 4570 1080
rect 10538 -16 11752 1078
<< viali >>
rect 3558 1893 3663 1959
rect 3746 1919 3812 1981
rect 3965 1900 4033 1999
rect 11047 1885 11181 1959
rect 11235 1919 11301 1985
rect 11454 1882 11540 2005
rect 3558 1285 3704 1333
rect 3752 1083 3818 1149
rect 10931 1062 10993 1132
rect 11207 1109 11273 1175
rect 11330 1112 11373 1241
rect 3921 910 4000 1023
rect 11597 843 11677 1035
<< metal1 >>
rect 2980 2904 4612 3038
rect 7527 2904 9159 3038
rect 10503 2904 11506 3038
rect 3537 2359 4017 2904
rect 11026 2361 11506 2904
rect 1979 2127 1989 2185
rect 2252 2127 2262 2185
rect 6543 2128 6553 2185
rect 6817 2128 6827 2185
rect 9526 2126 9536 2180
rect 9796 2126 9806 2180
rect 3959 1999 4039 2011
rect 11448 2005 11546 2017
rect 3734 1981 3824 1987
rect 3546 1959 3675 1965
rect 3546 1929 3558 1959
rect 3663 1929 3675 1959
rect 3538 1785 3548 1929
rect 3675 1785 3685 1929
rect 3734 1919 3746 1981
rect 3812 1919 3824 1981
rect 3734 1913 3824 1919
rect 3955 1900 3965 1999
rect 4033 1900 4043 1999
rect 11223 1985 11313 1991
rect 11035 1959 11193 1965
rect 3959 1888 4039 1900
rect 11035 1885 11047 1959
rect 11181 1885 11193 1959
rect 11223 1919 11235 1985
rect 11301 1919 11313 1985
rect 11223 1913 11313 1919
rect 11035 1879 11193 1885
rect 11444 1882 11454 2005
rect 11540 1882 11550 2005
rect 11448 1870 11546 1882
rect 2949 1370 4573 1698
rect 10503 1370 11694 1698
rect 3546 1333 3716 1339
rect 3546 1279 3558 1333
rect 3704 1279 3716 1333
rect 11324 1252 11379 1253
rect 11324 1241 11350 1252
rect 11195 1175 11285 1181
rect 3740 1149 3830 1155
rect 3740 1083 3752 1149
rect 3818 1083 3830 1149
rect 10925 1132 10999 1144
rect 3740 1077 3830 1083
rect 10901 1046 10911 1132
rect 10996 1046 11006 1132
rect 11195 1109 11207 1175
rect 11273 1109 11285 1175
rect 11195 1103 11285 1109
rect 11324 1112 11330 1241
rect 11421 1113 11431 1252
rect 11373 1112 11379 1113
rect 11324 1100 11379 1112
rect 11591 1038 11683 1047
rect 11591 1035 11727 1038
rect 3915 1023 4006 1035
rect 1969 888 1979 942
rect 2245 888 2255 942
rect 3911 910 3921 1023
rect 4000 910 4010 1023
rect 3915 898 4006 910
rect 6527 888 6537 941
rect 6850 888 6860 941
rect 9524 883 9534 937
rect 9798 883 9808 937
rect 11591 843 11597 1035
rect 11677 843 11727 1035
rect 11591 831 11683 843
rect 3537 164 4017 715
rect 11053 164 11533 736
rect 2959 30 4591 164
rect 7544 30 9176 164
rect 10496 30 11533 164
<< via1 >>
rect 1989 2127 2252 2185
rect 6553 2128 6817 2185
rect 9536 2126 9796 2180
rect 3548 1893 3558 1929
rect 3558 1893 3663 1929
rect 3663 1893 3675 1929
rect 3548 1785 3675 1893
rect 3746 1919 3812 1981
rect 3965 1900 4033 1999
rect 11047 1885 11181 1959
rect 11235 1919 11301 1985
rect 11454 1882 11540 2005
rect 3558 1285 3704 1333
rect 3558 1279 3704 1285
rect 11350 1241 11421 1252
rect 3752 1083 3818 1149
rect 10911 1062 10931 1132
rect 10931 1062 10993 1132
rect 10993 1062 10996 1132
rect 10911 1046 10996 1062
rect 11207 1109 11273 1175
rect 11350 1113 11373 1241
rect 11373 1113 11421 1241
rect 1979 888 2245 942
rect 3921 910 4000 1023
rect 6537 888 6850 941
rect 9534 883 9798 937
<< metal2 >>
rect 1989 2191 2256 2201
rect 1989 2117 2256 2127
rect 6548 2190 6820 2200
rect 6548 2111 6820 2121
rect 9528 2191 9800 2201
rect 9528 2111 9800 2121
rect 3060 2010 3812 2076
rect 2763 1597 2823 1607
rect 3060 1565 3126 2010
rect 3746 1981 3812 2010
rect 3548 1929 3675 1939
rect 3746 1909 3812 1919
rect 3965 1999 4033 2009
rect 11454 2005 11540 2015
rect 11235 1985 11301 1995
rect 11047 1959 11181 1969
rect 3675 1785 3676 1798
rect 3548 1775 3676 1785
rect 3549 1694 3676 1775
rect 2823 1499 3126 1565
rect 3256 1567 3676 1694
rect 2763 1459 2823 1469
rect 1970 943 2254 953
rect 1970 861 2254 871
rect 3256 -184 3383 1567
rect 3558 1333 3704 1343
rect 3558 1269 3704 1279
rect 3580 403 3640 1269
rect 3752 1150 3818 1159
rect 3965 1150 4033 1900
rect 10651 1888 11047 1954
rect 10317 1608 10377 1618
rect 4817 1573 4877 1583
rect 4263 1566 4817 1567
rect 3752 1149 4033 1150
rect 3818 1083 4033 1149
rect 3752 1082 4033 1083
rect 4226 1501 4817 1566
rect 3752 1073 3818 1082
rect 3921 1023 4000 1033
rect 4226 1004 4292 1501
rect 4817 1483 4877 1493
rect 10651 1580 10717 1888
rect 11047 1875 11181 1885
rect 11235 1715 11301 1919
rect 11454 1872 11540 1882
rect 10377 1514 10717 1580
rect 10773 1649 11301 1715
rect 10317 1470 10377 1480
rect 4000 938 4292 1004
rect 6537 950 6850 951
rect 6523 941 6876 950
rect 6523 940 6537 941
rect 6850 940 6876 941
rect 3921 900 4000 910
rect 6523 859 6876 869
rect 9523 946 9823 956
rect 9523 859 9823 869
rect 3559 393 3664 403
rect 3559 224 3664 234
rect 3580 -26 3640 224
rect 7123 -26 7183 810
rect 7800 476 7866 800
rect 10773 476 10839 1649
rect 11461 1539 11527 1872
rect 11207 1479 11527 1539
rect 11207 1175 11273 1479
rect 11350 1252 11421 1262
rect 10894 1140 11014 1150
rect 11207 1099 11273 1109
rect 11339 1113 11350 1248
rect 11339 1103 11421 1113
rect 10894 954 11014 964
rect 7800 410 10839 476
rect 11339 -26 11399 1103
rect 3580 -86 11399 -26
rect 3256 -196 11063 -184
rect 3256 -306 10863 -196
rect 11050 -306 11063 -196
rect 3256 -311 11063 -306
rect 10863 -316 11050 -311
<< via2 >>
rect 1989 2185 2256 2191
rect 1989 2127 2252 2185
rect 2252 2127 2256 2185
rect 6548 2185 6820 2190
rect 6548 2128 6553 2185
rect 6553 2128 6817 2185
rect 6817 2128 6820 2185
rect 6548 2121 6820 2128
rect 9528 2180 9800 2191
rect 9528 2126 9536 2180
rect 9536 2126 9796 2180
rect 9796 2126 9800 2180
rect 9528 2121 9800 2126
rect 2763 1469 2823 1597
rect 1970 942 2254 943
rect 1970 888 1979 942
rect 1979 888 2245 942
rect 2245 888 2254 942
rect 1970 871 2254 888
rect 4817 1493 4877 1573
rect 10317 1480 10377 1608
rect 6523 888 6537 940
rect 6537 888 6850 940
rect 6850 888 6876 940
rect 6523 869 6876 888
rect 9523 937 9823 946
rect 9523 883 9534 937
rect 9534 883 9798 937
rect 9798 883 9823 937
rect 9523 869 9823 883
rect 3559 234 3664 393
rect 10894 1132 11014 1140
rect 10894 1046 10911 1132
rect 10911 1046 10996 1132
rect 10996 1046 11014 1132
rect 10894 964 11014 1046
rect 10863 -306 11050 -196
<< metal3 >>
rect 247 804 307 2264
rect 1978 2123 1988 2199
rect 2270 2123 2280 2199
rect 6538 2190 6830 2195
rect 1979 2122 2266 2123
rect 6538 2121 6548 2190
rect 6820 2121 6830 2190
rect 6538 2116 6830 2121
rect 9486 2112 9496 2202
rect 9810 2112 9820 2202
rect 10307 1608 10387 1613
rect 2753 1597 2833 1602
rect 2753 1469 2763 1597
rect 2823 1469 2833 1597
rect 4807 1573 4887 1578
rect 4807 1493 4817 1573
rect 4877 1493 4887 1573
rect 7379 1504 7861 1564
rect 4807 1488 4887 1493
rect 10307 1480 10317 1608
rect 10377 1480 10387 1608
rect 10307 1475 10387 1480
rect 2753 1464 2833 1469
rect 10893 1145 11020 1154
rect 10884 1140 11024 1145
rect 10884 964 10894 1140
rect 11014 964 11024 1140
rect 10884 959 11024 964
rect 1951 861 1961 951
rect 2267 861 2277 951
rect 9513 946 9833 951
rect 6513 940 6886 945
rect 6513 869 6523 940
rect 6876 869 6886 940
rect 6513 864 6886 869
rect 9513 869 9523 946
rect 9823 869 9833 946
rect 9513 864 9833 869
rect 238 388 311 789
rect 3549 393 3674 398
rect 224 267 234 388
rect 311 267 321 388
rect 238 263 311 267
rect 3549 234 3559 393
rect 3664 234 3674 393
rect 3549 229 3674 234
rect 10893 -184 11020 959
rect 10892 -191 11020 -184
rect 10853 -196 11060 -191
rect 10853 -306 10863 -196
rect 11050 -306 11060 -196
rect 10853 -311 11060 -306
<< via3 >>
rect 1988 2191 2270 2199
rect 1988 2127 1989 2191
rect 1989 2127 2256 2191
rect 2256 2127 2270 2191
rect 1988 2123 2270 2127
rect 6548 2121 6820 2190
rect 9496 2191 9810 2202
rect 9496 2121 9528 2191
rect 9528 2121 9800 2191
rect 9800 2121 9810 2191
rect 9496 2112 9810 2121
rect 1961 943 2267 951
rect 1961 871 1970 943
rect 1970 871 2254 943
rect 2254 871 2267 943
rect 1961 861 2267 871
rect 6523 869 6876 940
rect 9523 869 9823 946
rect 234 267 311 388
rect 3559 234 3664 393
<< metal4 >>
rect 1983 2203 9735 2204
rect 1983 2202 9811 2203
rect 1983 2199 9496 2202
rect 1983 2123 1988 2199
rect 2270 2190 9496 2199
rect 2270 2123 6548 2190
rect 1983 2121 6548 2123
rect 6820 2121 9496 2190
rect 1983 2112 9496 2121
rect 9810 2112 9811 2202
rect 9495 2111 9811 2112
rect 1960 951 9783 952
rect 1960 861 1961 951
rect 2267 947 9783 951
rect 2267 946 9824 947
rect 2267 940 9523 946
rect 2267 869 6523 940
rect 6876 869 9523 940
rect 9823 869 9824 946
rect 2267 868 9824 869
rect 2267 861 9783 868
rect 1960 860 9783 861
rect 3558 393 3665 394
rect 233 388 312 389
rect 233 267 234 388
rect 311 377 312 388
rect 3558 377 3559 393
rect 311 267 3559 377
rect 233 266 312 267
rect 3558 234 3559 267
rect 3664 234 3665 393
rect 3558 233 3665 234
use sky130_fd_sc_hs__mux2_1  sky130_fd_sc_hs__mux2_1_0
timestamp 1623986409
transform 1 0 10830 0 -1 1419
box -38 -49 902 715
use sky130_fd_sc_hs__or2_1  sky130_fd_sc_hs__or2_1_0
timestamp 1624049879
transform 1 0 3537 0 1 1649
box -38 -49 518 715
use sky130_fd_sc_hs__or2_1  sky130_fd_sc_hs__or2_1_1
timestamp 1624049879
transform 1 0 11026 0 1 1649
box -38 -49 518 715
use sky130_fd_sc_hs__and2_1  sky130_fd_sc_hs__and2_1_0
timestamp 1624049879
transform 1 0 3537 0 -1 1419
box -38 -49 518 715
use DFlipFlop  DFlipFlop_0
timestamp 1624885207
transform 1 0 1244 0 1 0
box -1244 0 1740 3068
use DFlipFlop  DFlipFlop_1
timestamp 1624885207
transform 1 0 5814 0 1 0
box -1244 0 1740 3068
use DFlipFlop  DFlipFlop_2
timestamp 1624885207
transform 1 0 8798 0 -1 3068
box -1244 0 1740 3068
<< labels >>
rlabel metal4 2267 860 6523 952 1 CLK
rlabel metal4 2270 2112 6548 2204 1 nCLK
rlabel metal1 11677 843 11727 1038 1 CLK_23
rlabel metal1 2980 2904 4612 3038 1 vdd
rlabel metal1 2949 1370 4573 1698 1 vss
rlabel metal4 311 267 3559 377 1 nCLK_23
rlabel metal2 3256 -311 10863 -184 1 MC
rlabel metal2 3060 1499 3126 2076 1 Q1
rlabel metal3 7379 1504 7861 1564 1 Q2
rlabel metal2 10651 1888 11047 1954 1 Q2_d
<< end >>
