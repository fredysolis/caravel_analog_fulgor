magic
tech sky130A
magscale 1 2
timestamp 1624397222
<< nwell >>
rect 18234 4138 21604 4172
<< pwell >>
rect 21025 7249 22667 7283
rect 22739 7250 26841 7284
rect 26993 4400 27027 7051
rect 26993 1269 27027 3920
rect 21025 1046 22667 1080
rect 22739 1047 26841 1081
<< psubdiff >>
rect 21025 7249 21121 7283
rect 21767 7249 21925 7283
rect 22571 7249 22667 7283
rect 22739 7250 22835 7284
rect 26745 7250 26841 7284
rect 18334 5923 18358 7205
rect 20851 5923 20875 7205
rect 26993 6989 27027 7051
rect 26993 5221 27027 5379
rect 26993 4400 27027 4447
rect 26993 3873 27027 3920
rect 26993 2941 27027 3099
rect 18338 1138 18362 2420
rect 20855 1138 20879 2420
rect 26993 1269 27027 1331
rect 21025 1046 21121 1080
rect 21767 1046 21925 1080
rect 22571 1046 22667 1080
rect 22739 1047 22835 1081
rect 26745 1047 26841 1081
<< nsubdiff >>
rect 18234 4138 18330 4172
rect 19840 4138 19998 4172
rect 21508 4138 21604 4172
<< psubdiffcont >>
rect 21121 7249 21767 7283
rect 21925 7249 22571 7283
rect 22835 7250 26745 7284
rect 18358 5923 20851 7205
rect 26993 5379 27027 6989
rect 26993 4447 27027 5221
rect 26993 3099 27027 3873
rect 18362 1138 20855 2420
rect 26993 1331 27027 2941
rect 21121 1046 21767 1080
rect 21925 1046 22571 1080
rect 22835 1047 26745 1081
<< nsubdiffcont >>
rect 18330 4138 19840 4172
rect 19998 4138 21508 4172
<< locali >>
rect 18342 5923 18358 7205
rect 20851 5923 20867 7205
rect 18346 1138 18362 2420
rect 20855 1138 20871 2420
<< viali >>
rect 21025 7249 21121 7283
rect 21121 7249 21767 7283
rect 21767 7249 21925 7283
rect 21925 7249 22571 7283
rect 22571 7249 22667 7283
rect 22739 7250 22835 7284
rect 22835 7250 26745 7284
rect 26745 7250 26841 7284
rect 18358 5923 20851 7205
rect 26993 6989 27027 7051
rect 26993 5379 27027 6989
rect 26993 5221 27027 5379
rect 26993 4447 27027 5221
rect 26993 4400 27027 4447
rect 18234 4138 18330 4172
rect 18330 4138 19840 4172
rect 19840 4138 19998 4172
rect 19998 4138 21508 4172
rect 21508 4138 21604 4172
rect 26993 3873 27027 3920
rect 26993 3099 27027 3873
rect 26993 2941 27027 3099
rect 18362 1138 20855 2420
rect 26993 1331 27027 2941
rect 26993 1269 27027 1331
rect 21025 1046 21121 1080
rect 21121 1046 21767 1080
rect 21767 1046 21925 1080
rect 21925 1046 22571 1080
rect 22571 1046 22667 1080
rect 22739 1047 22835 1081
rect 22835 1047 26745 1081
rect 26745 1047 26841 1081
<< metal1 >>
rect -4991 11573 -4981 12019
rect -4333 11856 -4323 12019
rect -4333 11826 -198 11856
rect -4333 11743 -4273 11826
rect -301 11743 -198 11826
rect -4333 11721 -198 11743
rect 7413 11792 7708 11855
rect -4333 11573 -4323 11721
rect 7413 11692 7547 11792
rect 7674 11692 7708 11792
rect 7413 11639 7708 11692
rect 7298 10621 18864 10683
rect -3030 10141 -3020 10587
rect -2372 10515 -2362 10587
rect 7298 10552 9156 10621
rect -2372 10466 -188 10515
rect -2372 10231 -2293 10466
rect -318 10231 -188 10466
rect -2372 10187 -188 10231
rect 7298 10286 7940 10552
rect 8700 10289 9156 10552
rect 18767 10289 18864 10621
rect 8700 10286 18864 10289
rect 7298 10187 18864 10286
rect -2372 10141 -2362 10187
rect 18368 10108 18864 10187
rect -4967 8592 -4957 9038
rect -4309 8981 -4299 9038
rect -4309 8951 -210 8981
rect -4309 8684 -4173 8951
rect -505 8684 -210 8951
rect -4309 8653 -210 8684
rect 7023 8946 12143 8981
rect 7023 8842 9064 8946
rect 7023 8687 7537 8842
rect 7688 8687 9064 8842
rect -4309 8592 -4299 8653
rect 7023 8624 9064 8687
rect 11661 8910 12143 8946
rect 11661 8624 11766 8910
rect 12080 8624 12143 8910
rect 7023 8571 12143 8624
rect 6160 8096 14598 8113
rect 6160 7969 9070 8096
rect 14582 7969 14598 8096
rect 6160 7958 14598 7969
rect 14341 7920 14598 7958
rect 6398 7533 9126 7712
rect 6398 7531 9001 7533
rect -3020 7076 -3010 7522
rect -2362 7448 -2352 7522
rect 6674 7471 9001 7531
rect -2362 7399 -204 7448
rect -2362 7167 -2268 7399
rect -443 7167 -204 7399
rect -2362 7119 -204 7167
rect 6674 7205 7936 7471
rect 8696 7205 9001 7471
rect -2362 7076 -2352 7119
rect 6674 6953 9001 7205
rect 11249 6504 11259 6610
rect 11353 6504 11363 6610
rect -4970 5531 -4960 5977
rect -4312 5913 -4302 5977
rect -4312 5860 -89 5913
rect -4312 5630 -4206 5860
rect -493 5630 -89 5860
rect -4312 5585 -89 5630
rect 5819 5746 9205 5996
rect -4312 5531 -4302 5585
rect 5819 5562 7506 5746
rect 7708 5562 9205 5746
rect 5819 5437 9205 5562
rect 12670 5544 13227 7679
rect 14341 6257 14357 7920
rect 14579 6436 14598 7920
rect 18368 7462 18460 10108
rect 18773 7462 18864 10108
rect 18368 7211 18864 7462
rect 21025 7283 22739 7284
rect 22667 7282 22739 7283
rect 18346 7205 20863 7211
rect 14579 6341 15829 6436
rect 14579 6313 14598 6341
rect 14579 6257 14599 6313
rect 14341 6109 14599 6257
rect 14341 6056 14598 6109
rect -3024 4004 -3014 4450
rect -2366 4379 -2356 4450
rect -2366 4334 -195 4379
rect -2366 4102 -2293 4334
rect -311 4102 -195 4334
rect -2366 4051 -195 4102
rect -2366 4004 -2356 4051
rect -4955 1523 -4945 1969
rect -4297 1911 -4287 1969
rect -242 1911 170 2845
rect 7412 2673 7422 2892
rect 7737 2673 7747 2892
rect 13666 2667 13676 2699
rect -4297 1855 170 1911
rect -4297 1620 -4217 1855
rect -353 1620 170 1855
rect -4297 1583 170 1620
rect -4297 1523 -4287 1583
rect -242 1366 170 1583
rect -242 988 454 1366
rect 13603 1118 13676 2667
rect 13920 2667 13930 2699
rect 13920 1118 14010 2667
rect 14393 1971 14488 2240
rect 15734 1971 15829 6341
rect 18346 5923 18358 7205
rect 20851 5923 20863 7205
rect 21015 7093 21025 7282
rect 26841 7093 26851 7282
rect 21734 6516 21744 6620
rect 21940 6516 21950 6620
rect 18346 5917 20863 5923
rect 18976 5035 18986 5130
rect 19121 5035 19131 5130
rect 28363 6957 28373 7403
rect 29021 6957 29031 7403
rect 18236 4172 18246 4216
rect 18357 4172 18367 4216
rect 18453 4172 18463 4344
rect 18236 4105 18246 4138
rect 18357 4105 18367 4138
rect 18453 3979 18463 4138
rect 21653 3979 21663 4344
rect 21815 4035 21825 4290
rect 26610 4035 26620 4290
rect 26993 3920 27027 4400
rect 18975 3197 18985 3292
rect 19120 3197 19130 3292
rect 14393 1876 15829 1971
rect 18350 2420 20867 2426
rect 13603 1094 14010 1118
rect 18197 1463 18201 1512
rect 18197 1094 18206 1463
rect 18350 1138 18362 2420
rect 20855 1138 20867 2420
rect 21735 1699 21745 1803
rect 21941 1699 21951 1803
rect 27070 3749 27075 4585
rect 18350 1132 20867 1138
rect 12803 895 12813 1085
rect 13201 895 13211 1085
rect 13603 954 18979 1094
rect 21015 1046 21025 1235
rect 26841 1046 26851 1235
rect 13603 168 13721 954
rect 12256 132 13721 168
rect 18694 132 18979 954
rect 12256 28 18979 132
<< via1 >>
rect -4981 11573 -4333 12019
rect -4273 11743 -301 11826
rect 7547 11692 7674 11792
rect -3020 10141 -2372 10587
rect -2293 10231 -318 10466
rect 7940 10286 8700 10552
rect 9156 10289 18767 10621
rect -4957 8592 -4309 9038
rect -4173 8684 -505 8951
rect 7537 8687 7688 8842
rect 9064 8624 11661 8946
rect 11766 8624 12080 8910
rect 9070 7969 14582 8096
rect -3010 7076 -2362 7522
rect -2268 7167 -443 7399
rect 7936 7205 8696 7471
rect 11259 6504 11353 6610
rect -4960 5531 -4312 5977
rect -4206 5630 -493 5860
rect 7506 5562 7708 5746
rect 14357 6257 14579 7920
rect 18460 7462 18773 10108
rect -3014 4004 -2366 4450
rect -2293 4102 -311 4334
rect -4945 1523 -4297 1969
rect 7422 2673 7737 2892
rect -4217 1620 -353 1855
rect 13676 1118 13920 2699
rect 18358 5923 20851 7205
rect 21025 7249 22667 7282
rect 22667 7250 22739 7282
rect 22739 7250 26841 7282
rect 22667 7249 26841 7250
rect 21025 7093 26841 7249
rect 21744 6516 21940 6620
rect 18986 5035 19121 5130
rect 28373 6957 29021 7403
rect 18246 4172 18357 4216
rect 18463 4172 21653 4344
rect 18246 4138 18357 4172
rect 18463 4138 21604 4172
rect 21604 4138 21653 4172
rect 18246 4105 18357 4138
rect 18463 3979 21653 4138
rect 21825 4035 26610 4290
rect 18985 3197 19120 3292
rect 18362 1138 20855 2420
rect 21745 1699 21941 1803
rect 12813 895 13201 1085
rect 21025 1081 26841 1235
rect 21025 1080 22739 1081
rect 21025 1046 22667 1080
rect 22667 1047 22739 1080
rect 22739 1047 26841 1081
rect 22667 1046 26841 1047
rect 13721 132 18694 954
<< metal2 >>
rect -4981 12019 -4333 12029
rect -4333 11836 -4249 11840
rect -4333 11826 -301 11836
rect -4333 11743 -4273 11826
rect -4333 11733 -301 11743
rect 7547 11792 7674 11802
rect -4333 11730 -4249 11733
rect -4981 11563 -4333 11573
rect 7547 11560 7674 11692
rect -3020 10587 -2372 10597
rect -2372 10476 -2217 10489
rect -2372 10466 -318 10476
rect -2372 10231 -2293 10466
rect -2372 10221 -318 10231
rect -2372 10200 -2217 10221
rect -3020 10131 -2372 10141
rect -4957 9038 -4309 9048
rect -4309 8961 -4120 8962
rect -4309 8951 -505 8961
rect -4309 8684 -4173 8951
rect 7548 8852 7672 11560
rect 9156 10621 18767 10631
rect 7940 10552 8700 10562
rect 7940 10276 8700 10286
rect 9156 10279 18767 10289
rect 18460 10108 18773 10118
rect 9064 8946 11661 8956
rect -4309 8674 -505 8684
rect 7537 8842 7688 8852
rect 7537 8677 7688 8687
rect -4309 8673 -4120 8674
rect -4957 8582 -4309 8592
rect -3010 7522 -2362 7532
rect -2268 7399 -443 7409
rect -2268 7157 -443 7167
rect -3010 7066 -2362 7076
rect 5620 6412 6084 6624
rect -4960 5977 -4312 5987
rect -4312 5870 -4159 5884
rect -4312 5860 -493 5870
rect -4312 5630 -4206 5860
rect -4312 5620 -493 5630
rect -4312 5595 -4159 5620
rect -4960 5521 -4312 5531
rect -3014 4450 -2366 4460
rect -2366 4344 -2194 4361
rect -2366 4334 -311 4344
rect -2366 4102 -2293 4334
rect -2366 4092 -311 4102
rect -2366 4072 -2194 4092
rect -3014 3994 -2366 4004
rect 5873 3175 6083 6412
rect 7548 5756 7672 8677
rect 9064 8614 11661 8624
rect 11766 8910 12080 8920
rect 11766 8614 12080 8624
rect 9070 8096 14582 8106
rect 9070 7959 14582 7969
rect 14357 7920 14579 7930
rect 7936 7471 8696 7481
rect 7936 7195 8696 7205
rect 11259 6610 11353 6620
rect 11259 6494 11353 6504
rect 19819 8935 20467 8945
rect 19819 8479 20467 8489
rect 18460 7452 18773 7462
rect 19830 7215 20449 8479
rect 28373 7403 29021 7413
rect 21025 7282 28373 7292
rect 14357 6247 14579 6257
rect 18358 7205 20851 7215
rect 26841 7093 28373 7282
rect 21025 7083 28373 7093
rect 28373 6947 29021 6957
rect 21744 6620 21940 6630
rect 21744 6506 21940 6516
rect 18358 5913 20851 5923
rect 7506 5746 7708 5756
rect 7506 5552 7708 5562
rect -117 2965 6083 3175
rect -4945 1969 -4297 1979
rect -4297 1865 -4118 1889
rect -4297 1855 -353 1865
rect -4297 1620 -4217 1855
rect -4297 1610 -353 1620
rect -4297 1600 -4118 1610
rect -4945 1513 -4297 1523
rect -117 579 93 2965
rect 7548 2902 7672 5552
rect 27126 5401 27326 5411
rect 15141 5204 15341 5214
rect 26993 5194 27027 5401
rect 27126 5184 27326 5194
rect 18986 5130 19121 5140
rect 18986 5025 19121 5035
rect 15141 4681 15341 4691
rect 30366 4380 31014 4390
rect 18463 4344 21653 4354
rect 8505 4334 8631 4344
rect 8505 4256 8631 4266
rect 18246 4216 18357 4226
rect 15465 4105 18246 4216
rect 18246 4095 18357 4105
rect 8505 4046 8631 4056
rect 8505 3968 8631 3978
rect 21825 4290 30366 4300
rect 26610 4035 30366 4290
rect 21825 4025 30366 4035
rect 26541 4021 30366 4025
rect 18463 3969 21653 3979
rect 30366 3924 31014 3934
rect 15141 3621 15341 3631
rect 18985 3292 19120 3302
rect 18985 3187 19120 3197
rect 27126 3126 27326 3136
rect 15141 3098 15341 3108
rect 26993 2919 27027 3126
rect 27126 2909 27326 2919
rect 7422 2892 7737 2902
rect 7422 2663 7737 2673
rect 13676 2699 13920 2709
rect 2703 2553 2856 2563
rect 2703 2463 2856 2473
rect 9277 2471 9430 2481
rect 9277 2381 9430 2391
rect -117 500 -107 579
rect 77 500 93 579
rect -117 480 93 500
rect 239 2280 380 2365
rect 239 2270 409 2280
rect -3006 419 -2358 429
rect 239 341 380 2270
rect 18362 2420 20855 2430
rect 21745 1803 21941 1813
rect 21745 1689 21941 1699
rect 28405 1367 29053 1377
rect 18362 1128 20855 1138
rect 21025 1235 28405 1245
rect 13676 1108 13920 1118
rect 12813 1085 13201 1095
rect 12813 885 13201 895
rect 13721 954 18694 964
rect -2358 65 380 341
rect 13721 122 18694 132
rect 239 40 380 65
rect -3006 -37 -2358 -27
rect 19830 -155 20449 1128
rect 26841 1046 28405 1235
rect 21025 1036 28405 1046
rect 28405 911 29053 921
rect 19819 -165 20467 -155
rect 19819 -621 20467 -611
<< via2 >>
rect -4981 11573 -4333 12019
rect -3020 10141 -2372 10587
rect -4957 8592 -4309 9038
rect 7940 10286 8700 10552
rect -3010 7076 -2362 7522
rect -4960 5531 -4312 5977
rect -3014 4004 -2366 4450
rect 11766 8624 12080 8910
rect 7936 7205 8696 7471
rect 11259 6504 11353 6610
rect 19819 8489 20467 8935
rect 28373 6957 29021 7403
rect 21744 6516 21940 6620
rect -4945 1523 -4297 1969
rect 15141 4691 15341 5204
rect 27126 5194 27326 5401
rect 8505 4266 8631 4334
rect 8505 3978 8631 4046
rect 30366 3934 31014 4380
rect 15141 3108 15341 3621
rect 27126 2919 27326 3126
rect 2703 2473 2856 2553
rect 9277 2391 9430 2471
rect -107 500 77 579
rect -3006 -27 -2358 419
rect 21745 1699 21941 1803
rect 12813 895 13201 1085
rect 15257 783 15796 949
rect 28405 921 29053 1367
rect 19819 -611 20467 -165
<< metal3 >>
rect -4991 12019 -4323 12024
rect -4991 11573 -4981 12019
rect -4333 11573 -4323 12019
rect -4991 11568 -4323 11573
rect -3030 10587 -2362 10592
rect -3030 10141 -3020 10587
rect -2372 10141 -2362 10587
rect -3030 10136 -2362 10141
rect 7797 10552 8854 12355
rect 7797 10286 7940 10552
rect 8700 10286 8854 10552
rect -4967 9038 -4299 9043
rect -4967 8592 -4957 9038
rect -4309 8592 -4299 9038
rect -4967 8587 -4299 8592
rect -3020 7522 -2352 7527
rect -3020 7076 -3010 7522
rect -2362 7076 -2352 7522
rect -3020 7071 -2352 7076
rect -4970 5977 -4302 5982
rect -4970 5531 -4960 5977
rect -4312 5531 -4302 5977
rect -4970 5526 -4302 5531
rect -709 4799 -603 9765
rect 7797 7471 8854 10286
rect 19809 8935 20477 8940
rect 11756 8910 12090 8915
rect 11756 8624 11766 8910
rect 12081 8625 12091 8910
rect 12080 8624 12090 8625
rect 11756 8619 12090 8624
rect 11766 8605 12080 8619
rect 19809 8489 19819 8935
rect 20467 8489 20477 8935
rect 19809 8484 20477 8489
rect 7797 7205 7936 7471
rect 8696 7205 8854 7471
rect 7797 4525 8854 7205
rect 28363 7403 29031 7408
rect 10855 6954 10865 7060
rect 10959 6954 10969 7060
rect 11459 6958 11469 7064
rect 11563 6958 11573 7064
rect 12458 6951 12468 7057
rect 12562 6951 12572 7057
rect 28363 6957 28373 7403
rect 29021 6957 29031 7403
rect 28363 6952 29031 6957
rect 21734 6620 21950 6625
rect 11249 6610 11363 6615
rect 11249 6504 11259 6610
rect 11353 6504 11363 6610
rect 11249 6499 11363 6504
rect 14157 6163 15942 6545
rect 21734 6516 21744 6620
rect 21940 6516 21950 6620
rect 21734 6511 21950 6516
rect 15131 5204 15351 5209
rect 15131 4691 15141 5204
rect 15341 4691 15351 5204
rect 15131 4686 15351 4691
rect -3024 4450 -2356 4455
rect -3024 4004 -3014 4450
rect -2366 4004 -2356 4450
rect 8495 4334 8641 4339
rect 8495 4266 8505 4334
rect 8631 4266 8641 4334
rect 8495 4261 8641 4266
rect -3024 3999 -2356 4004
rect 8495 4046 8641 4051
rect 8495 3978 8505 4046
rect 8631 3978 8641 4046
rect 8495 3973 8641 3978
rect 15131 3621 15351 3626
rect 15131 3108 15141 3621
rect 15341 3108 15351 3621
rect 15131 3103 15351 3108
rect 2693 2553 2866 2558
rect 2693 2473 2703 2553
rect 2856 2473 2866 2553
rect 6820 2486 6830 2566
rect 6983 2486 6993 2566
rect 2693 2468 2866 2473
rect 9267 2471 9440 2476
rect 9267 2391 9277 2471
rect 9430 2391 9440 2471
rect 9267 2386 9440 2391
rect 15560 2115 15942 6163
rect 17802 5620 17812 5768
rect 18033 5620 18043 5768
rect 27116 5401 27336 5406
rect 27116 5194 27126 5401
rect 27326 5194 27336 5401
rect 27116 5189 27336 5194
rect 30356 4380 31024 4385
rect 30356 3934 30366 4380
rect 31014 3934 31024 4380
rect 30356 3929 31024 3934
rect 27116 3126 27336 3131
rect 27116 2919 27126 3126
rect 27326 2919 27336 3126
rect 27116 2914 27336 2919
rect 17802 2552 17812 2700
rect 18033 2552 18043 2700
rect -4955 1969 -4287 1974
rect -4955 1523 -4945 1969
rect -4297 1523 -4287 1969
rect 14152 1733 15942 2115
rect 21735 1803 21951 1808
rect -4955 1518 -4287 1523
rect 12803 1085 13211 1090
rect 12803 895 12813 1085
rect 13201 895 13211 1085
rect 15316 954 15765 1733
rect 21735 1699 21745 1803
rect 21941 1699 21951 1803
rect 21735 1694 21951 1699
rect 28395 1367 29063 1372
rect 12803 890 13211 895
rect 15247 949 15806 954
rect 15247 783 15257 949
rect 15796 783 15806 949
rect 28395 921 28405 1367
rect 29053 921 29063 1367
rect 28395 916 29063 921
rect 15247 778 15806 783
rect -117 579 87 584
rect -117 500 -107 579
rect 77 574 87 579
rect 77 512 200 574
rect 77 500 87 512
rect -117 495 87 500
rect -3016 419 -2348 424
rect -3016 -27 -3006 419
rect -2358 -27 -2348 419
rect -3016 -32 -2348 -27
rect 19809 -165 20477 -160
rect 19809 -611 19819 -165
rect 20467 -611 20477 -165
rect 19809 -616 20477 -611
<< via3 >>
rect -4981 11573 -4333 12019
rect -3020 10141 -2372 10587
rect -4957 8592 -4309 9038
rect -3010 7076 -2362 7522
rect -4960 5531 -4312 5977
rect 11766 8625 12080 8910
rect 12080 8625 12081 8910
rect 19819 8489 20467 8935
rect 10865 6954 10959 7060
rect 11469 6958 11563 7064
rect 12468 6951 12562 7057
rect 28373 6957 29021 7403
rect 11259 6504 11353 6610
rect 15141 4691 15341 5204
rect -3014 4004 -2366 4450
rect 8505 4266 8631 4334
rect 8505 3978 8631 4046
rect 15141 3108 15341 3621
rect 2703 2473 2856 2553
rect 6830 2486 6983 2566
rect 9277 2391 9430 2471
rect 17812 5620 18033 5768
rect 27126 5194 27326 5401
rect 30366 3934 31014 4380
rect 27126 2919 27326 3126
rect 17812 2552 18033 2700
rect -4945 1523 -4297 1969
rect 12813 895 13201 1085
rect 28405 921 29053 1367
rect -3006 -27 -2358 419
rect 19819 -611 20467 -165
<< metal4 >>
rect -4982 12019 -4332 12020
rect -4982 11573 -4981 12019
rect -4333 11573 -4332 12019
rect -4982 11572 -4332 11573
rect -3021 10587 -2371 10588
rect -3021 10141 -3020 10587
rect -2372 10141 -2371 10587
rect -3021 10140 -2371 10141
rect -4958 9038 -4308 9039
rect -4958 8592 -4957 9038
rect -4309 8592 -4308 9038
rect -4958 8591 -4308 8592
rect -3011 7522 -2361 7523
rect -3011 7076 -3010 7522
rect -2362 7076 -2361 7522
rect -3011 7075 -2361 7076
rect -4961 5977 -4311 5978
rect -4961 5531 -4960 5977
rect -4312 5531 -4311 5977
rect -4961 5530 -4311 5531
rect -3015 4450 -2365 4451
rect -3015 4004 -3014 4450
rect -2366 4004 -2365 4450
rect -3015 4003 -2365 4004
rect -1112 3556 -968 11010
rect 8025 4047 8152 12638
rect 8505 4339 8632 12638
rect 11710 9974 30894 9975
rect 11710 9532 30333 9974
rect 11710 8910 12153 9532
rect 11710 8625 11766 8910
rect 12081 8625 12153 8910
rect 11468 7064 11564 7065
rect 10864 7060 10960 7061
rect 10864 6954 10865 7060
rect 10959 6954 10960 7060
rect 11468 6958 11469 7064
rect 11563 6958 11564 7064
rect 11468 6957 11564 6958
rect 10864 6953 10960 6954
rect 11258 6610 11354 6611
rect 11258 6504 11259 6610
rect 11353 6504 11354 6610
rect 11258 6503 11354 6504
rect 11710 5473 12153 8625
rect 19818 8935 20468 8936
rect 19818 8489 19819 8935
rect 20467 8489 20468 8935
rect 19818 8488 20468 8489
rect 28372 7403 29022 7404
rect 12467 7057 12563 7058
rect 12467 6951 12468 7057
rect 12562 6951 12563 7057
rect 28372 6957 28373 7403
rect 29021 6957 29022 7403
rect 28372 6956 29022 6957
rect 12467 6950 12563 6951
rect 17640 5768 18034 5769
rect 17640 5620 17812 5768
rect 18033 5620 18034 5768
rect 17640 5619 18034 5620
rect 17640 5205 17840 5619
rect 15140 5204 17840 5205
rect 15140 4691 15141 5204
rect 15341 5005 17840 5204
rect 27125 5401 27327 5402
rect 27125 5194 27126 5401
rect 27326 5194 27327 5401
rect 27125 5193 27327 5194
rect 15341 4691 15342 5005
rect 15140 4690 15342 4691
rect 8504 4334 8632 4339
rect 8504 4266 8505 4334
rect 8631 4266 8632 4334
rect 8504 4265 8632 4266
rect 30365 4380 31015 4381
rect 8025 4046 8632 4047
rect 8025 3978 8505 4046
rect 8631 3978 8632 4046
rect 8025 3977 8632 3978
rect 30365 3934 30366 4380
rect 31014 3934 31015 4380
rect 30365 3933 31015 3934
rect 15140 3621 15342 3622
rect 15140 3108 15141 3621
rect 15341 3307 15342 3621
rect 15341 3108 17841 3307
rect 15140 3107 17841 3108
rect 17641 2701 17841 3107
rect 27125 3126 27327 3127
rect 27125 2919 27126 3126
rect 27326 2919 27327 3126
rect 27125 2918 27327 2919
rect 17641 2700 18034 2701
rect 6829 2566 6984 2567
rect 2702 2553 2857 2554
rect 2702 2473 2703 2553
rect 2856 2473 2857 2553
rect 6829 2486 6830 2566
rect 6983 2486 6984 2566
rect 17641 2552 17812 2700
rect 18033 2552 18034 2700
rect 17641 2551 18034 2552
rect 6829 2485 6984 2486
rect 2702 2472 2857 2473
rect 9276 2471 9431 2472
rect 9276 2391 9277 2471
rect 9430 2391 9431 2471
rect 9276 2390 9431 2391
rect -4946 1969 -4296 1970
rect -4946 1523 -4945 1969
rect -4297 1523 -4296 1969
rect -4946 1522 -4296 1523
rect 28404 1367 29054 1368
rect 12812 1085 13202 1086
rect 12812 993 12813 1085
rect 12799 895 12813 993
rect 13201 993 13202 1085
rect 13201 895 13242 993
rect 28404 921 28405 1367
rect 29053 921 29054 1367
rect 28404 920 29054 921
rect -3007 419 -2357 420
rect -3007 -27 -3006 419
rect -2358 -27 -2357 419
rect -3007 -28 -2357 -27
rect 12799 -503 13242 895
rect -4286 -946 13242 -503
rect 19818 -165 20468 -164
rect 19818 -611 19819 -165
rect 20467 -611 20468 -165
rect 19818 -612 20468 -611
<< via4 >>
rect -4981 11573 -4333 12019
rect -3020 10141 -2372 10587
rect -4957 8592 -4309 9038
rect -3010 7076 -2362 7522
rect -4960 5531 -4312 5977
rect -3014 4004 -2366 4450
rect 30333 9528 30981 9974
rect 19819 8489 20467 8935
rect 28373 6957 29021 7403
rect 30366 3934 31014 4380
rect -4945 1523 -4297 1969
rect 28405 921 29053 1367
rect -3006 -27 -2358 419
rect -4934 -948 -4286 -502
rect 19819 -611 20467 -165
<< metal5 >>
rect -4855 12043 -4412 12726
rect -5005 12019 -4309 12043
rect -5005 11573 -4981 12019
rect -4333 11573 -4309 12019
rect -5005 11549 -4309 11573
rect -4855 9062 -4412 11549
rect -2910 10611 -2467 12726
rect -3044 10587 -2348 10611
rect -3044 10141 -3020 10587
rect -2372 10141 -2348 10587
rect -3044 10117 -2348 10141
rect -4981 9038 -4285 9062
rect -4981 8592 -4957 9038
rect -4309 8592 -4285 9038
rect -4981 8568 -4285 8592
rect -4855 6001 -4412 8568
rect -2910 7546 -2467 10117
rect 19795 8935 20491 8959
rect 19795 8489 19819 8935
rect 20467 8929 20491 8935
rect 28506 8929 28949 12726
rect 30451 9998 30894 12726
rect 30309 9974 31005 9998
rect 30309 9528 30333 9974
rect 30981 9528 31005 9974
rect 30309 9504 31005 9528
rect 20467 8489 28949 8929
rect 19795 8486 28949 8489
rect 19795 8465 20491 8486
rect -3034 7522 -2338 7546
rect -3034 7076 -3010 7522
rect -2362 7076 -2338 7522
rect 28506 7427 28949 8486
rect -3034 7052 -2338 7076
rect 28349 7403 29045 7427
rect -4984 5977 -4288 6001
rect -4984 5531 -4960 5977
rect -4312 5531 -4288 5977
rect -4984 5507 -4288 5531
rect -4855 1993 -4412 5507
rect -2910 4474 -2467 7052
rect 28349 6957 28373 7403
rect 29021 6957 29045 7403
rect 28349 6933 29045 6957
rect -3038 4450 -2342 4474
rect -3038 4004 -3014 4450
rect -2366 4004 -2342 4450
rect -3038 3980 -2342 4004
rect -4969 1969 -4273 1993
rect -4969 1523 -4945 1969
rect -4297 1523 -4273 1969
rect -4969 1499 -4273 1523
rect -4855 -478 -4412 1499
rect -2910 443 -2467 3980
rect 28506 1391 28949 6933
rect 30451 4404 30894 9504
rect 30342 4380 31038 4404
rect 30342 3934 30366 4380
rect 31014 3934 31038 4380
rect 30342 3910 31038 3934
rect 28381 1367 29077 1391
rect 28381 921 28405 1367
rect 29053 921 29077 1367
rect 28381 897 29077 921
rect -3030 419 -2334 443
rect -3030 -27 -3006 419
rect -2358 -27 -2334 419
rect -3030 -51 -2334 -27
rect -2910 -129 -2467 -51
rect 19795 -162 20491 -141
rect 28506 -162 28949 897
rect 30451 -147 30894 3910
rect 19795 -165 28949 -162
rect -4958 -502 -4262 -478
rect -4958 -948 -4934 -502
rect -4286 -948 -4262 -502
rect 19795 -611 19819 -165
rect 20467 -605 28949 -165
rect 20467 -611 20491 -605
rect 19795 -635 20491 -611
rect -4958 -972 -4262 -948
use source_follower_buff_diff  source_follower_buff_diff_0
timestamp 1624113565
transform 1 0 17170 0 1 1168
box 863 -174 10692 6158
use res_amp_sync_v2  res_amp_sync_v2_0
timestamp 1624397222
transform 1 0 -899 0 1 4870
box -92 -2189 8342 7015
use res_amp_lin_prog  res_amp_lin_prog_0
timestamp 1624397222
transform 1 0 -5726 0 1 -7077
box 5835 7077 21302 14799
<< labels >>
rlabel metal4 8534 12559 8597 12604 1 inn
rlabel metal4 8060 12573 8123 12618 1 inp
rlabel metal4 -1064 10918 -1018 10975 1 clkn
rlabel space -742 9560 -696 9617 1 clkp
rlabel metal4 27211 5274 27257 5331 1 outp
rlabel metal4 27221 2994 27267 3051 1 outn
rlabel metal4 2733 2487 2790 2523 1 delay_reg2
rlabel metal4 9327 2414 9384 2450 1 delay_reg0
rlabel metal4 6829 2485 6886 2521 1 delay_reg1
rlabel metal4 10864 6953 10960 7061 1 iref_reg0
rlabel metal4 11468 6957 11564 7065 1 iref_reg1
rlabel metal4 12467 6950 12563 7058 1 iref_reg2
rlabel metal5 -2784 12535 -2629 12632 1 avss1p8
rlabel metal5 -4717 12539 -4562 12636 1 avdd1p8
rlabel metal4 11259 6504 11353 6610 1 iref0
rlabel via1 18986 5035 19121 5130 1 iref1
rlabel via1 18985 3197 19120 3292 1 iref3
rlabel metal3 21744 6516 21940 6620 1 iref2
rlabel metal3 21745 1699 21941 1803 1 iref4
<< end >>
