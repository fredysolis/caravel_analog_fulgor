magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< pwell >>
rect -257 -327 257 327
<< nmos >>
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
<< ndiff >>
rect -221 288 -159 300
rect -221 -288 -209 288
rect -175 -288 -159 288
rect -221 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 221 300
rect 159 -288 175 288
rect 209 -288 221 288
rect 159 -300 221 -288
<< ndiffc >>
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
<< poly >>
rect -257 326 257 499
rect -159 300 -129 326
rect -63 300 -33 326
rect 33 300 63 326
rect 129 300 159 326
rect -159 -322 -129 -300
rect -63 -322 -33 -300
rect 33 -322 63 -300
rect 129 -322 159 -300
rect -257 -404 257 -322
<< locali >>
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
<< viali >>
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
<< metal1 >>
rect -257 353 257 435
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -343 -169 -288
rect -119 288 -73 353
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -343 23 -288
rect 73 288 119 353
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -343 215 -288
rect -257 -425 257 -343
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -306 -457 306 457
string parameters w 3 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
