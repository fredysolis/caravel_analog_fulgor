magic
tech sky130A
magscale 1 2
timestamp 1624020278
<< metal3 >>
rect -4309 50 -141 4250
rect 10 4222 4309 4250
rect 10 78 4225 4222
rect 4289 78 4309 4222
rect 10 50 4309 78
rect -4309 -4250 -141 -50
rect 10 -78 4309 -50
rect 10 -4222 4225 -78
rect 4289 -4222 4309 -78
rect 10 -4250 4309 -4222
<< via3 >>
rect 4225 78 4289 4222
rect 4225 -4222 4289 -78
<< mimcap >>
rect -4209 4110 -209 4150
rect -4209 190 -4169 4110
rect -249 190 -209 4110
rect -4209 150 -209 190
rect 110 4110 4110 4150
rect 110 190 150 4110
rect 4070 190 4110 4110
rect 110 150 4110 190
rect -4209 -190 -209 -150
rect -4209 -4110 -4169 -190
rect -249 -4110 -209 -190
rect -4209 -4150 -209 -4110
rect 110 -190 4110 -150
rect 110 -4110 150 -190
rect 4070 -4110 4110 -190
rect 110 -4150 4110 -4110
<< mimcapcontact >>
rect -4169 190 -249 4110
rect 150 190 4070 4110
rect -4169 -4110 -249 -190
rect 150 -4110 4070 -190
<< metal4 >>
rect -2261 4111 -2157 4300
rect 2058 4111 2162 4300
rect 4178 4238 4282 4300
rect 4178 4222 4305 4238
rect -4170 4110 -248 4111
rect -4170 190 -4169 4110
rect -249 190 -248 4110
rect -4170 189 -248 190
rect 149 4110 4071 4111
rect 149 190 150 4110
rect 4070 190 4071 4110
rect 149 189 4071 190
rect -2261 -189 -2157 189
rect 2058 -189 2162 189
rect 4178 78 4225 4222
rect 4289 78 4305 4222
rect 4178 62 4305 78
rect 4178 -62 4282 62
rect 4178 -78 4305 -62
rect -4170 -190 -248 -189
rect -4170 -4110 -4169 -190
rect -249 -4110 -248 -190
rect -4170 -4111 -248 -4110
rect 149 -190 4071 -189
rect 149 -4110 150 -190
rect 4070 -4110 4071 -190
rect 149 -4111 4071 -4110
rect -2261 -4300 -2157 -4111
rect 2058 -4300 2162 -4111
rect 4178 -4222 4225 -78
rect 4289 -4222 4305 -78
rect 4178 -4238 4305 -4222
rect 4178 -4300 4282 -4238
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 10 50 4210 4250
string parameters w 20 l 20 val 815.2 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
