magic
tech sky130A
magscale 1 2
timestamp 1624653480
<< poly >>
rect 420 -552 654 -486
rect 588 -670 654 -552
rect 588 -736 833 -670
<< metal1 >>
rect -11 -76 1267 2
rect 198 -670 290 -580
rect 332 -760 424 -670
rect -11 -1360 1267 -1282
<< metal2 >>
rect 586 -424 678 -131
rect 616 -583 1041 -517
rect 616 -679 682 -583
rect 404 -745 682 -679
rect 41 -1224 111 -929
rect 1145 -1225 1215 -930
use trans_gate_mux2to8  trans_gate_mux2to8_1
timestamp 1624653480
transform -1 0 1203 0 -1 -723
box -64 -725 579 637
use trans_gate_mux2to8  trans_gate_mux2to8_0
timestamp 1624653480
transform 1 0 53 0 -1 -723
box -64 -725 579 637
<< labels >>
rlabel metal2 586 -424 678 -131 1 in_a
rlabel metal1 -11 -76 1267 2 1 vss
rlabel metal1 -11 -1360 1267 -1282 1 vdd
rlabel metal2 41 -1224 111 -929 1 out_a_0
rlabel metal2 1145 -1225 1215 -930 1 out_a_1
rlabel metal1 198 -670 290 -580 1 select_0_neg
rlabel metal1 332 -760 424 -670 1 select_0
<< end >>
