magic
tech sky130A
magscale 1 2
timestamp 1624046389
<< nwell >>
rect -935 -303 935 303
<< pmos >>
rect -735 -84 -705 84
rect -639 -84 -609 84
rect -543 -84 -513 84
rect -447 -84 -417 84
rect -351 -84 -321 84
rect -255 -84 -225 84
rect -159 -84 -129 84
rect -63 -84 -33 84
rect 33 -84 63 84
rect 129 -84 159 84
rect 225 -84 255 84
rect 321 -84 351 84
rect 417 -84 447 84
rect 513 -84 543 84
rect 609 -84 639 84
rect 705 -84 735 84
<< pdiff >>
rect -797 72 -735 84
rect -797 -72 -785 72
rect -751 -72 -735 72
rect -797 -84 -735 -72
rect -705 72 -639 84
rect -705 -72 -689 72
rect -655 -72 -639 72
rect -705 -84 -639 -72
rect -609 72 -543 84
rect -609 -72 -593 72
rect -559 -72 -543 72
rect -609 -84 -543 -72
rect -513 72 -447 84
rect -513 -72 -497 72
rect -463 -72 -447 72
rect -513 -84 -447 -72
rect -417 72 -351 84
rect -417 -72 -401 72
rect -367 -72 -351 72
rect -417 -84 -351 -72
rect -321 72 -255 84
rect -321 -72 -305 72
rect -271 -72 -255 72
rect -321 -84 -255 -72
rect -225 72 -159 84
rect -225 -72 -209 72
rect -175 -72 -159 72
rect -225 -84 -159 -72
rect -129 72 -63 84
rect -129 -72 -113 72
rect -79 -72 -63 72
rect -129 -84 -63 -72
rect -33 72 33 84
rect -33 -72 -17 72
rect 17 -72 33 72
rect -33 -84 33 -72
rect 63 72 129 84
rect 63 -72 79 72
rect 113 -72 129 72
rect 63 -84 129 -72
rect 159 72 225 84
rect 159 -72 175 72
rect 209 -72 225 72
rect 159 -84 225 -72
rect 255 72 321 84
rect 255 -72 271 72
rect 305 -72 321 72
rect 255 -84 321 -72
rect 351 72 417 84
rect 351 -72 367 72
rect 401 -72 417 72
rect 351 -84 417 -72
rect 447 72 513 84
rect 447 -72 463 72
rect 497 -72 513 72
rect 447 -84 513 -72
rect 543 72 609 84
rect 543 -72 559 72
rect 593 -72 609 72
rect 543 -84 609 -72
rect 639 72 705 84
rect 639 -72 655 72
rect 689 -72 705 72
rect 639 -84 705 -72
rect 735 72 797 84
rect 735 -72 751 72
rect 785 -72 797 72
rect 735 -84 797 -72
<< pdiffc >>
rect -785 -72 -751 72
rect -689 -72 -655 72
rect -593 -72 -559 72
rect -497 -72 -463 72
rect -401 -72 -367 72
rect -305 -72 -271 72
rect -209 -72 -175 72
rect -113 -72 -79 72
rect -17 -72 17 72
rect 79 -72 113 72
rect 175 -72 209 72
rect 271 -72 305 72
rect 367 -72 401 72
rect 463 -72 497 72
rect 559 -72 593 72
rect 655 -72 689 72
rect 751 -72 785 72
<< nsubdiff >>
rect -899 233 -803 267
rect 803 233 899 267
rect -899 171 -865 233
rect 865 171 899 233
rect -899 -267 -865 -171
rect 865 -267 899 -171
<< nsubdiffcont >>
rect -803 233 803 267
rect -899 -171 -865 171
rect 865 -171 899 171
<< poly >>
rect -752 110 753 181
rect -735 84 -705 110
rect -639 84 -609 110
rect -543 84 -513 110
rect -447 84 -417 110
rect -351 84 -321 110
rect -255 84 -225 110
rect -159 84 -129 110
rect -63 84 -33 110
rect 33 84 63 110
rect 129 84 159 110
rect 225 84 255 110
rect 321 84 351 110
rect 417 84 447 110
rect 513 84 543 110
rect 609 84 639 110
rect 705 84 735 110
rect -735 -110 -705 -84
rect -639 -110 -609 -84
rect -543 -110 -513 -84
rect -447 -110 -417 -84
rect -351 -110 -321 -84
rect -255 -110 -225 -84
rect -159 -110 -129 -84
rect -63 -110 -33 -84
rect 33 -110 63 -84
rect 129 -110 159 -84
rect 225 -110 255 -84
rect 321 -110 351 -84
rect 417 -110 447 -84
rect 513 -110 543 -84
rect 609 -110 639 -84
rect 705 -110 735 -84
rect -753 -181 752 -110
<< locali >>
rect -899 233 -803 267
rect 803 233 899 267
rect -899 171 -865 233
rect 865 171 899 233
rect -785 72 -751 88
rect -785 -88 -751 -72
rect -689 72 -655 88
rect -689 -88 -655 -72
rect -593 72 -559 88
rect -593 -88 -559 -72
rect -497 72 -463 88
rect -497 -88 -463 -72
rect -401 72 -367 88
rect -401 -88 -367 -72
rect -305 72 -271 88
rect -305 -88 -271 -72
rect -209 72 -175 88
rect -209 -88 -175 -72
rect -113 72 -79 88
rect -113 -88 -79 -72
rect -17 72 17 88
rect -17 -88 17 -72
rect 79 72 113 88
rect 79 -88 113 -72
rect 175 72 209 88
rect 175 -88 209 -72
rect 271 72 305 88
rect 271 -88 305 -72
rect 367 72 401 88
rect 367 -88 401 -72
rect 463 72 497 88
rect 463 -88 497 -72
rect 559 72 593 88
rect 559 -88 593 -72
rect 655 72 689 88
rect 655 -88 689 -72
rect 751 72 785 88
rect 751 -88 785 -72
rect -899 -267 -865 -171
rect 865 -267 899 -171
<< viali >>
rect -785 -72 -751 72
rect -689 -72 -655 72
rect -593 -72 -559 72
rect -497 -72 -463 72
rect -401 -72 -367 72
rect -305 -72 -271 72
rect -209 -72 -175 72
rect -113 -72 -79 72
rect -17 -72 17 72
rect 79 -72 113 72
rect 175 -72 209 72
rect 271 -72 305 72
rect 367 -72 401 72
rect 463 -72 497 72
rect 559 -72 593 72
rect 655 -72 689 72
rect 751 -72 785 72
<< metal1 >>
rect -791 72 -745 84
rect -791 -72 -785 72
rect -751 -72 -745 72
rect -791 -84 -745 -72
rect -695 72 -649 84
rect -695 -72 -689 72
rect -655 -72 -649 72
rect -695 -84 -649 -72
rect -599 72 -553 84
rect -599 -72 -593 72
rect -559 -72 -553 72
rect -599 -84 -553 -72
rect -503 72 -457 84
rect -503 -72 -497 72
rect -463 -72 -457 72
rect -503 -84 -457 -72
rect -407 72 -361 84
rect -407 -72 -401 72
rect -367 -72 -361 72
rect -407 -84 -361 -72
rect -311 72 -265 84
rect -311 -72 -305 72
rect -271 -72 -265 72
rect -311 -84 -265 -72
rect -215 72 -169 84
rect -215 -72 -209 72
rect -175 -72 -169 72
rect -215 -84 -169 -72
rect -119 72 -73 84
rect -119 -72 -113 72
rect -79 -72 -73 72
rect -119 -84 -73 -72
rect -23 72 23 84
rect -23 -72 -17 72
rect 17 -72 23 72
rect -23 -84 23 -72
rect 73 72 119 84
rect 73 -72 79 72
rect 113 -72 119 72
rect 73 -84 119 -72
rect 169 72 215 84
rect 169 -72 175 72
rect 209 -72 215 72
rect 169 -84 215 -72
rect 265 72 311 84
rect 265 -72 271 72
rect 305 -72 311 72
rect 265 -84 311 -72
rect 361 72 407 84
rect 361 -72 367 72
rect 401 -72 407 72
rect 361 -84 407 -72
rect 457 72 503 84
rect 457 -72 463 72
rect 497 -72 503 72
rect 457 -84 503 -72
rect 553 72 599 84
rect 553 -72 559 72
rect 593 -72 599 72
rect 553 -84 599 -72
rect 649 72 695 84
rect 649 -72 655 72
rect 689 -72 695 72
rect 649 -84 695 -72
rect 745 72 791 84
rect 745 -72 751 72
rect 785 -72 791 72
rect 745 -84 791 -72
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -882 -250 882 250
string parameters w 0.84 l 0.15 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
