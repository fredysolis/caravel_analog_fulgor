magic
tech sky130A
magscale 1 2
timestamp 1624046389
<< pwell >>
rect -935 -252 935 252
<< nmos >>
rect -735 -42 -705 42
rect -639 -42 -609 42
rect -543 -42 -513 42
rect -447 -42 -417 42
rect -351 -42 -321 42
rect -255 -42 -225 42
rect -159 -42 -129 42
rect -63 -42 -33 42
rect 33 -42 63 42
rect 129 -42 159 42
rect 225 -42 255 42
rect 321 -42 351 42
rect 417 -42 447 42
rect 513 -42 543 42
rect 609 -42 639 42
rect 705 -42 735 42
<< ndiff >>
rect -797 30 -735 42
rect -797 -30 -785 30
rect -751 -30 -735 30
rect -797 -42 -735 -30
rect -705 30 -639 42
rect -705 -30 -689 30
rect -655 -30 -639 30
rect -705 -42 -639 -30
rect -609 30 -543 42
rect -609 -30 -593 30
rect -559 -30 -543 30
rect -609 -42 -543 -30
rect -513 30 -447 42
rect -513 -30 -497 30
rect -463 -30 -447 30
rect -513 -42 -447 -30
rect -417 30 -351 42
rect -417 -30 -401 30
rect -367 -30 -351 30
rect -417 -42 -351 -30
rect -321 30 -255 42
rect -321 -30 -305 30
rect -271 -30 -255 30
rect -321 -42 -255 -30
rect -225 30 -159 42
rect -225 -30 -209 30
rect -175 -30 -159 30
rect -225 -42 -159 -30
rect -129 30 -63 42
rect -129 -30 -113 30
rect -79 -30 -63 30
rect -129 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 129 42
rect 63 -30 79 30
rect 113 -30 129 30
rect 63 -42 129 -30
rect 159 30 225 42
rect 159 -30 175 30
rect 209 -30 225 30
rect 159 -42 225 -30
rect 255 30 321 42
rect 255 -30 271 30
rect 305 -30 321 30
rect 255 -42 321 -30
rect 351 30 417 42
rect 351 -30 367 30
rect 401 -30 417 30
rect 351 -42 417 -30
rect 447 30 513 42
rect 447 -30 463 30
rect 497 -30 513 30
rect 447 -42 513 -30
rect 543 30 609 42
rect 543 -30 559 30
rect 593 -30 609 30
rect 543 -42 609 -30
rect 639 30 705 42
rect 639 -30 655 30
rect 689 -30 705 30
rect 639 -42 705 -30
rect 735 30 797 42
rect 735 -30 751 30
rect 785 -30 797 30
rect 735 -42 797 -30
<< ndiffc >>
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
<< psubdiff >>
rect -899 120 -865 216
rect 865 120 899 216
rect -899 -182 -865 -120
rect 865 -182 899 -120
rect -899 -216 -803 -182
rect 803 -216 899 -182
<< psubdiffcont >>
rect -899 -120 -865 120
rect 865 -120 899 120
rect -803 -216 803 -182
<< poly >>
rect -757 64 753 130
rect -735 42 -705 64
rect -639 42 -609 64
rect -543 42 -513 64
rect -447 42 -417 64
rect -351 42 -321 64
rect -255 42 -225 64
rect -159 42 -129 64
rect -63 42 -33 64
rect 33 42 63 64
rect 129 42 159 64
rect 225 42 255 64
rect 321 42 351 64
rect 417 42 447 64
rect 513 42 543 64
rect 609 42 639 64
rect 705 42 735 64
rect -735 -64 -705 -42
rect -639 -64 -609 -42
rect -543 -64 -513 -42
rect -447 -64 -417 -42
rect -351 -64 -321 -42
rect -255 -64 -225 -42
rect -159 -64 -129 -42
rect -63 -64 -33 -42
rect 33 -64 63 -42
rect 129 -64 159 -42
rect 225 -64 255 -42
rect 321 -64 351 -42
rect 417 -64 447 -42
rect 513 -64 543 -42
rect 609 -64 639 -42
rect 705 -64 735 -42
rect -753 -130 757 -64
<< locali >>
rect -899 120 -865 216
rect 865 120 899 216
rect -785 30 -751 46
rect -785 -46 -751 -30
rect -689 30 -655 46
rect -689 -46 -655 -30
rect -593 30 -559 46
rect -593 -46 -559 -30
rect -497 30 -463 46
rect -497 -46 -463 -30
rect -401 30 -367 46
rect -401 -46 -367 -30
rect -305 30 -271 46
rect -305 -46 -271 -30
rect -209 30 -175 46
rect -209 -46 -175 -30
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect 271 30 305 46
rect 271 -46 305 -30
rect 367 30 401 46
rect 367 -46 401 -30
rect 463 30 497 46
rect 463 -46 497 -30
rect 559 30 593 46
rect 559 -46 593 -30
rect 655 30 689 46
rect 655 -46 689 -30
rect 751 30 785 46
rect 751 -46 785 -30
rect -899 -182 -865 -120
rect 865 -182 899 -120
rect -899 -216 -803 -182
rect 803 -216 899 -182
<< viali >>
rect -785 -30 -751 30
rect -689 -30 -655 30
rect -593 -30 -559 30
rect -497 -30 -463 30
rect -401 -30 -367 30
rect -305 -30 -271 30
rect -209 -30 -175 30
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
rect 175 -30 209 30
rect 271 -30 305 30
rect 367 -30 401 30
rect 463 -30 497 30
rect 559 -30 593 30
rect 655 -30 689 30
rect 751 -30 785 30
<< metal1 >>
rect -791 30 -745 42
rect -791 -30 -785 30
rect -751 -30 -745 30
rect -791 -42 -745 -30
rect -695 30 -649 42
rect -695 -30 -689 30
rect -655 -30 -649 30
rect -695 -42 -649 -30
rect -599 30 -553 42
rect -599 -30 -593 30
rect -559 -30 -553 30
rect -599 -42 -553 -30
rect -503 30 -457 42
rect -503 -30 -497 30
rect -463 -30 -457 30
rect -503 -42 -457 -30
rect -407 30 -361 42
rect -407 -30 -401 30
rect -367 -30 -361 30
rect -407 -42 -361 -30
rect -311 30 -265 42
rect -311 -30 -305 30
rect -271 -30 -265 30
rect -311 -42 -265 -30
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect 265 30 311 42
rect 265 -30 271 30
rect 305 -30 311 30
rect 265 -42 311 -30
rect 361 30 407 42
rect 361 -30 367 30
rect 401 -30 407 30
rect 361 -42 407 -30
rect 457 30 503 42
rect 457 -30 463 30
rect 497 -30 503 30
rect 457 -42 503 -30
rect 553 30 599 42
rect 553 -30 559 30
rect 593 -30 599 30
rect 553 -42 599 -30
rect 649 30 695 42
rect 649 -30 655 30
rect 689 -30 695 30
rect 649 -42 695 -30
rect 745 30 791 42
rect 745 -30 751 30
rect 785 -30 791 30
rect 745 -42 791 -30
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -882 -199 882 199
string parameters w 0.420 l 0.150 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
