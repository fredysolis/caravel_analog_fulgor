magic
tech sky130A
magscale 1 2
timestamp 1624653480
<< nwell >>
rect -53 635 569 723
rect -53 -53 569 -47
<< pwell >>
rect -53 -64 569 -53
rect -53 -811 569 -723
<< psubdiff >>
rect 55 -775 79 -741
rect 437 -775 461 -741
<< nsubdiff >>
rect 55 653 79 687
rect 437 653 461 687
<< psubdiffcont >>
rect 79 -775 437 -741
<< nsubdiffcont >>
rect 79 653 437 687
<< poly >>
rect 147 69 371 135
rect 279 31 371 69
rect 279 -37 291 31
rect 359 -37 371 31
rect 279 -53 371 -37
rect 145 -69 237 -53
rect 145 -137 157 -69
rect 225 -137 237 -69
rect 145 -171 237 -137
rect 145 -237 369 -171
<< polycont >>
rect 291 -37 359 31
rect 157 -137 225 -69
<< locali >>
rect 279 31 371 47
rect 279 -37 291 31
rect 359 -37 371 31
rect 279 -53 371 -37
rect 145 -69 237 -53
rect 145 -137 157 -69
rect 225 -137 237 -69
rect 145 -153 237 -137
<< viali >>
rect -17 653 79 687
rect 79 653 437 687
rect 437 653 533 687
rect -17 565 533 599
rect 291 -37 359 31
rect 157 -137 225 -69
rect -17 -687 533 -653
rect -17 -775 79 -741
rect 79 -775 437 -741
rect 437 -775 533 -741
<< metal1 >>
rect -53 687 569 693
rect -53 653 -17 687
rect 533 653 569 687
rect -53 599 165 653
rect 217 599 569 653
rect -53 565 -17 599
rect 533 565 569 599
rect -53 559 165 565
rect 217 559 569 565
rect 45 462 329 508
rect 45 404 137 462
rect 283 404 329 462
rect 45 -171 97 404
rect 425 183 477 416
rect 187 120 233 178
rect 419 120 477 183
rect 187 74 477 120
rect 279 -53 291 37
rect 359 -53 371 37
rect 145 -143 157 -53
rect 225 -143 237 -53
rect 45 -217 329 -171
rect 45 -341 97 -217
rect 283 -263 329 -217
rect 45 -513 91 -341
rect 419 -343 477 74
rect 425 -455 477 -343
rect 419 -501 477 -455
rect 187 -559 233 -513
rect 379 -559 477 -501
rect 187 -605 477 -559
rect -53 -653 569 -647
rect -53 -687 -17 -653
rect 533 -687 569 -653
rect -53 -741 299 -687
rect 351 -741 569 -687
rect -53 -775 -17 -741
rect 533 -775 569 -741
rect -53 -781 569 -775
<< via1 >>
rect 165 653 217 663
rect 165 599 217 653
rect 165 565 217 599
rect 165 559 217 565
rect 291 31 359 37
rect 291 -37 359 31
rect 291 -53 359 -37
rect 157 -69 225 -53
rect 157 -137 225 -69
rect 157 -143 225 -137
rect 299 -687 351 -653
rect 299 -741 351 -687
rect 299 -757 351 -741
<< metal2 >>
rect 157 663 225 673
rect 157 559 165 663
rect 217 559 225 663
rect 157 -53 225 559
rect 157 -153 225 -143
rect 291 37 359 47
rect 291 -653 359 -53
rect 291 -757 299 -653
rect 351 -757 359 -653
rect 291 -766 359 -757
rect 299 -767 351 -766
use sky130_fd_pr__pfet_01v8_4798MH  sky130_fd_pr__pfet_01v8_4798MH_0
timestamp 1624062693
transform 1 0 258 0 1 291
box -311 -338 311 344
use sky130_fd_pr__nfet_01v8_BHR94T  sky130_fd_pr__nfet_01v8_BHR94T_0
timestamp 1624062693
transform 1 0 258 0 1 -388
box -311 -335 311 324
<< labels >>
rlabel metal1 217 599 569 653 1 vdd
rlabel metal1 -53 -741 299 -687 1 vss
rlabel space 419 -605 477 416 1 out
rlabel space 45 -513 97 508 1 in
<< end >>
