magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect 0 1216 918 1304
rect 0 598 96 1216
<< pwell >>
rect 0 0 918 88
<< psubdiff >>
rect 108 36 132 70
rect 786 36 810 70
<< nsubdiff >>
rect 204 1234 228 1268
rect 786 1234 810 1268
rect 36 1146 213 1180
rect 552 1146 616 1180
rect 36 1087 70 1146
rect 36 671 70 733
<< psubdiffcont >>
rect 132 36 786 70
<< nsubdiffcont >>
rect 228 1234 786 1268
rect 36 733 70 1087
<< poly >>
rect 170 720 326 786
rect 170 707 230 720
rect 170 625 183 707
rect 217 625 230 707
rect 392 669 458 786
rect 170 414 230 625
rect 296 609 458 669
rect 656 640 722 786
rect 296 584 356 609
rect 296 502 309 584
rect 343 502 356 584
rect 296 456 356 502
rect 656 558 667 640
rect 701 558 722 640
rect 656 410 722 558
<< polycont >>
rect 183 625 217 707
rect 309 502 343 584
rect 667 558 701 640
<< locali >>
rect 36 1087 70 1146
rect 36 671 70 733
rect 183 707 217 723
rect 183 609 217 625
rect 667 640 701 656
rect 309 584 343 600
rect 667 542 701 558
rect 309 486 343 502
<< viali >>
rect 36 1234 228 1268
rect 228 1234 786 1268
rect 786 1234 882 1268
rect 36 1146 882 1180
rect 183 625 217 707
rect 309 502 343 584
rect 667 558 701 640
rect 848 158 882 528
rect 36 124 882 158
rect 36 36 132 70
rect 132 36 786 70
rect 786 36 882 70
<< metal1 >>
rect 0 1268 918 1274
rect 0 1234 36 1268
rect 882 1234 918 1268
rect 0 1180 918 1234
rect 0 1146 36 1180
rect 882 1146 918 1180
rect 0 1140 918 1146
rect 240 997 286 1140
rect 432 985 478 1140
rect 640 988 686 1140
rect 336 789 382 829
rect 336 743 478 789
rect 177 707 223 719
rect 177 699 183 707
rect 36 633 183 699
rect 177 625 183 633
rect 217 625 223 707
rect 177 613 223 625
rect 432 631 478 743
rect 661 640 707 652
rect 661 631 667 640
rect 303 584 349 596
rect 303 576 309 584
rect 36 510 309 576
rect 303 502 309 510
rect 343 502 349 584
rect 303 490 349 502
rect 432 565 667 631
rect 432 462 478 565
rect 661 558 667 565
rect 701 558 707 640
rect 661 546 707 558
rect 336 416 478 462
rect 336 388 382 416
rect 144 164 190 307
rect 528 164 574 308
rect 640 164 686 302
rect 766 298 812 997
rect 842 528 888 540
rect 842 164 848 528
rect 0 158 848 164
rect 882 164 888 528
rect 0 124 36 158
rect 882 124 918 164
rect 0 70 918 124
rect 0 36 36 70
rect 882 36 918 70
rect 0 30 918 36
rect 884 28 918 30
use sky130_fd_pr__pfet_01v8_7T83YG  sky130_fd_pr__pfet_01v8_7T83YG_0
timestamp 1624049879
transform 1 0 359 0 1 907
box -263 -309 263 309
use sky130_fd_pr__nfet_01v8_ZCYAJJ  sky130_fd_pr__nfet_01v8_ZCYAJJ_0
timestamp 1624049879
transform 1 0 359 0 1 343
box -359 -255 359 255
use sky130_fd_pr__nfet_01v8_ZXAV3F  sky130_fd_pr__nfet_01v8_ZXAV3F_0
timestamp 1624049879
transform 1 0 707 0 1 343
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_4F7GBC  sky130_fd_pr__pfet_01v8_4F7GBC_0
timestamp 1624049879
transform 1 0 707 0 1 907
box -211 -309 211 309
<< labels >>
rlabel metal1 0 70 918 124 1 vss
rlabel metal1 0 1180 918 1234 1 vdd
rlabel metal1 36 633 183 699 1 A
rlabel metal1 36 510 309 576 1 B
rlabel metal1 766 298 812 997 1 out
<< end >>
