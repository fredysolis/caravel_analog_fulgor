magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect 2872 706 3790 1304
rect 3241 700 3768 706
<< metal1 >>
rect 1390 1234 1400 1268
rect 0 1180 1400 1234
rect 1390 1146 1400 1180
rect 1472 1234 1482 1268
rect 2836 1234 3504 1274
rect 1472 1180 3504 1234
rect 1472 1146 1482 1180
rect 2836 1140 3504 1180
rect 0 652 210 718
rect 3150 676 3504 1140
rect 3754 97 3775 101
rect 2123 36 2176 39
rect 175 30 2786 36
rect 0 -30 2872 30
rect 2952 -26 2962 78
rect 3014 -26 3024 78
rect 3651 45 3661 97
rect 3765 45 3775 97
rect 3754 35 3775 45
rect 175 -36 2123 -30
rect 2159 -36 2786 -30
rect 3752 -32 3775 -22
rect 2865 -164 2919 -58
rect 3651 -84 3661 -32
rect 3765 -84 3775 -32
rect 3716 -88 3775 -84
rect 2872 -434 2919 -164
rect 0 -718 210 -652
rect 1390 -1180 1400 -1146
rect 0 -1234 1400 -1180
rect 1390 -1268 1400 -1234
rect 1472 -1180 1482 -1146
rect 1472 -1234 2872 -1180
rect 1472 -1268 1482 -1234
<< via1 >>
rect 1400 1146 1472 1268
rect 2962 -26 3014 78
rect 3661 45 3765 97
rect 3661 -84 3765 -32
rect 1400 -1268 1472 -1146
<< metal2 >>
rect 1400 1268 1472 1278
rect 1400 1136 1472 1146
rect 2802 572 3790 624
rect 2159 36 2211 436
rect 3686 107 3738 572
rect 3661 97 3765 107
rect 2962 78 3014 88
rect 2159 -26 2962 36
rect 3014 -26 3024 36
rect 3661 35 3765 45
rect 2159 -36 3024 -26
rect 3661 -32 3765 -22
rect 2159 -436 2211 -36
rect 3661 -94 3765 -84
rect 3686 -572 3738 -94
rect 2806 -624 3789 -572
rect 1400 -1146 1472 -1136
rect 1400 -1278 1472 -1268
<< via2 >>
rect 1400 1146 1472 1268
rect 1400 -1268 1472 -1146
<< metal3 >>
rect 1390 1268 1482 1273
rect 1390 1146 1400 1268
rect 1472 1146 1482 1268
rect 1390 1141 1482 1146
rect 1400 -1141 1472 1141
rect 1390 -1146 1482 -1141
rect 1390 -1268 1400 -1146
rect 1472 -1268 1482 -1146
rect 1390 -1273 1482 -1268
use dff_pfd  dff_pfd_1
timestamp 1624049879
transform 1 0 0 0 -1 0
box 0 0 2872 1304
use dff_pfd  dff_pfd_0
timestamp 1624049879
transform 1 0 0 0 1 0
box 0 0 2872 1304
use and_pfd  and_pfd_0
timestamp 1624049879
transform -1 0 3790 0 1 -598
box 0 0 918 1304
<< labels >>
rlabel metal1 0 652 210 718 1 A
rlabel metal1 0 -718 210 -652 1 B
rlabel metal1 0 -30 2872 30 1 vss
rlabel metal2 2802 572 3790 624 1 Up
rlabel metal2 2806 -624 3789 -572 1 Down
rlabel metal1 0 1180 3504 1234 1 vdd
rlabel metal2 2159 -436 2211 436 1 Reset
<< end >>
