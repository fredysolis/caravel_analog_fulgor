magic
tech sky130A
magscale 1 2
timestamp 1623248172
<< nwell >>
rect -363 1865 931 1954
rect -363 1858 911 1865
rect -363 1835 -280 1858
<< pwell >>
rect 500 321 931 387
rect 922 -121 931 321
rect 500 -193 931 -121
rect 924 -226 931 -193
rect -354 -904 929 -869
rect -363 -1001 929 -904
rect -363 -1002 -231 -1001
rect 799 -1002 929 -1001
<< psubdiff >>
rect 608 -174 632 -140
rect 790 -174 814 -140
rect -255 -966 -231 -932
rect 799 -966 823 -932
<< nsubdiff >>
rect -255 1884 -231 1918
rect 799 1884 823 1918
<< psubdiffcont >>
rect 632 -174 790 -140
rect -231 -966 799 -932
<< nsubdiffcont >>
rect -231 1884 799 1918
<< viali >>
rect -327 1884 -231 1918
rect -231 1884 799 1918
rect 799 1884 895 1918
rect -327 1795 895 1829
rect -327 1197 -293 1795
rect 861 1197 895 1795
rect -327 1163 895 1197
rect 536 -85 886 -51
rect 536 -174 632 -140
rect 632 -174 790 -140
rect 790 -174 886 -140
rect -327 -263 895 -229
rect -327 -843 -293 -263
rect 861 -843 895 -263
rect -327 -877 895 -843
rect -327 -966 -231 -932
rect -231 -966 799 -932
rect 799 -966 895 -932
<< metal1 >>
rect -363 1918 931 1924
rect -363 1884 -327 1918
rect 895 1884 931 1918
rect -363 1829 931 1884
rect -363 1163 -327 1829
rect -293 1789 861 1795
rect -293 1203 -287 1789
rect -180 1693 -170 1745
rect 738 1693 748 1745
rect -126 1636 -73 1646
rect -219 1203 -173 1348
rect -126 1346 -73 1356
rect 65 1636 119 1646
rect 65 1356 66 1636
rect 257 1637 311 1646
rect -27 1203 19 1351
rect 65 1346 119 1356
rect 165 1203 211 1358
rect 310 1357 311 1637
rect 450 1636 502 1646
rect 257 1346 311 1357
rect 357 1203 403 1360
rect 642 1636 694 1646
rect 450 1346 502 1356
rect 549 1203 595 1360
rect 642 1346 694 1356
rect 741 1203 787 1359
rect 855 1203 861 1789
rect -293 1197 861 1203
rect 895 1163 931 1829
rect -363 1157 931 1163
rect 68 1108 500 1157
rect 209 897 261 907
rect 209 607 261 617
rect 68 361 78 413
rect 286 361 296 413
rect 356 361 366 413
rect 490 361 500 413
rect 631 361 641 413
rect 693 361 703 413
rect 209 167 261 177
rect 644 173 690 361
rect 772 89 818 556
rect 209 27 261 37
rect 619 8 629 60
rect 733 8 743 60
rect 500 -51 931 -45
rect 500 -85 536 -51
rect 886 -85 931 -51
rect 500 -140 805 -85
rect 861 -140 931 -85
rect 500 -174 536 -140
rect 886 -174 931 -140
rect 68 -223 931 -174
rect -363 -229 931 -223
rect -363 -877 -327 -229
rect -293 -269 861 -263
rect -293 -837 -287 -269
rect -219 -403 -173 -269
rect -126 -413 -73 -403
rect -27 -404 19 -269
rect 165 -403 211 -269
rect 357 -403 403 -269
rect 549 -403 595 -269
rect 741 -403 787 -269
rect -126 -703 -73 -693
rect 65 -413 119 -403
rect 65 -693 66 -413
rect 65 -703 119 -693
rect 257 -412 311 -403
rect 310 -692 311 -412
rect 257 -703 311 -692
rect 450 -413 502 -403
rect 450 -703 502 -693
rect 642 -413 694 -403
rect 642 -703 694 -693
rect -180 -793 -170 -741
rect 738 -793 748 -741
rect 855 -837 861 -269
rect -293 -843 861 -837
rect 895 -877 931 -229
rect -363 -932 931 -877
rect -363 -966 -327 -932
rect 895 -966 931 -932
rect -363 -972 931 -966
<< via1 >>
rect -170 1693 738 1745
rect -126 1356 -73 1636
rect 66 1356 119 1636
rect 257 1357 310 1637
rect 450 1356 502 1636
rect 642 1356 694 1636
rect 209 617 261 897
rect 78 361 286 413
rect 366 361 490 413
rect 641 361 693 413
rect 209 37 261 167
rect 629 8 733 60
rect 805 -140 861 -85
rect 805 -141 861 -140
rect -126 -693 -73 -413
rect 66 -693 119 -413
rect 257 -692 310 -412
rect 450 -693 502 -413
rect 642 -693 694 -413
rect -170 -793 738 -741
<< metal2 >>
rect -180 1745 748 1755
rect -180 1693 -170 1745
rect 738 1693 748 1745
rect -180 1683 748 1693
rect -126 1636 -73 1646
rect 66 1636 119 1646
rect -73 1436 66 1563
rect -126 1346 -73 1356
rect 257 1637 310 1647
rect 119 1436 257 1563
rect 66 1346 119 1356
rect 209 1357 257 1436
rect 450 1636 502 1646
rect 310 1436 450 1563
rect 209 1347 310 1357
rect 642 1636 694 1646
rect 502 1436 642 1563
rect 209 897 261 1347
rect 450 1346 502 1356
rect 642 1346 694 1356
rect 639 1042 719 1046
rect 831 1042 851 1046
rect 209 607 261 617
rect 78 413 286 423
rect 68 361 78 413
rect 78 351 286 361
rect 366 413 490 423
rect 641 413 693 423
rect 490 361 641 413
rect 693 361 931 413
rect 366 351 490 361
rect 641 351 693 361
rect 209 167 261 177
rect 209 -402 261 37
rect 629 62 733 72
rect 629 -4 733 6
rect 805 -85 861 -75
rect 805 -151 861 -141
rect -126 -413 -73 -403
rect 66 -413 119 -403
rect -73 -613 66 -486
rect -126 -703 -73 -693
rect 209 -412 310 -402
rect 209 -486 257 -412
rect 119 -613 257 -486
rect 66 -703 119 -693
rect 450 -413 502 -403
rect 310 -613 450 -486
rect 257 -702 310 -692
rect 642 -413 694 -403
rect 502 -613 642 -486
rect 450 -703 502 -693
rect 642 -703 694 -693
rect -180 -741 748 -731
rect -180 -793 -170 -741
rect 738 -793 748 -741
rect -180 -802 748 -793
rect -180 -803 738 -802
<< via2 >>
rect 719 990 831 1046
rect 629 60 733 62
rect 629 8 733 60
rect 629 6 733 8
rect 805 -141 861 -85
<< metal3 >>
rect 709 1046 863 1051
rect 709 990 719 1046
rect 831 990 863 1046
rect 709 985 863 990
rect 619 62 743 67
rect 619 6 629 62
rect 733 6 743 62
rect 619 1 743 6
rect 650 -194 710 1
rect 803 -80 863 985
rect 795 -85 871 -80
rect 795 -141 805 -85
rect 861 -141 871 -85
rect 795 -146 871 -141
use cap_vco  cap_vco_0
timestamp 1623247475
transform 1 0 5 0 1 528
box 554 -6 926 514
use inverter_csvco  inverter_csvco_0
timestamp 1623162837
transform 1 0 68 0 1 387
box 0 -597 432 757
use sky130_fd_pr__pfet_01v8_8DL6ZL  sky130_fd_pr__pfet_01v8_8DL6ZL_0
timestamp 1622843784
transform -1 0 284 0 -1 1496
box -647 -369 647 369
use sky130_fd_pr__nfet_01v8_7H8F5S  sky130_fd_pr__nfet_01v8_7H8F5S_0
timestamp 1622843784
transform 1 0 284 0 -1 -553
box -647 -360 647 360
use sky130_fd_pr__nfet_01v8_EDT3AT  sky130_fd_pr__nfet_01v8_EDT3AT_0
timestamp 1623244079
transform 1 0 711 0 1 100
box -211 -221 211 221
<< labels >>
rlabel metal1 -363 1829 931 1884 1 vdd
rlabel metal1 -363 -932 931 -877 1 vss
rlabel metal2 -180 -803 -170 -731 1 vctrl
rlabel metal2 -180 1683 -170 1755 1 vbp
rlabel metal2 68 361 78 413 1 in
rlabel metal3 650 -194 710 6 1 D0
rlabel metal2 693 361 931 413 1 out
<< end >>
