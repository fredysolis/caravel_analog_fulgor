magic
tech sky130A
magscale 1 2
timestamp 1623985751
<< error_p >>
rect -1901 381 -1843 387
rect -1709 381 -1651 387
rect -1517 381 -1459 387
rect -1325 381 -1267 387
rect -1133 381 -1075 387
rect -941 381 -883 387
rect -749 381 -691 387
rect -557 381 -499 387
rect -365 381 -307 387
rect -173 381 -115 387
rect 19 381 77 387
rect 211 381 269 387
rect 403 381 461 387
rect 595 381 653 387
rect 787 381 845 387
rect 979 381 1037 387
rect 1171 381 1229 387
rect 1363 381 1421 387
rect 1555 381 1613 387
rect 1747 381 1805 387
rect -1901 347 -1889 381
rect -1709 347 -1697 381
rect -1517 347 -1505 381
rect -1325 347 -1313 381
rect -1133 347 -1121 381
rect -941 347 -929 381
rect -749 347 -737 381
rect -557 347 -545 381
rect -365 347 -353 381
rect -173 347 -161 381
rect 19 347 31 381
rect 211 347 223 381
rect 403 347 415 381
rect 595 347 607 381
rect 787 347 799 381
rect 979 347 991 381
rect 1171 347 1183 381
rect 1363 347 1375 381
rect 1555 347 1567 381
rect 1747 347 1759 381
rect -1901 341 -1843 347
rect -1709 341 -1651 347
rect -1517 341 -1459 347
rect -1325 341 -1267 347
rect -1133 341 -1075 347
rect -941 341 -883 347
rect -749 341 -691 347
rect -557 341 -499 347
rect -365 341 -307 347
rect -173 341 -115 347
rect 19 341 77 347
rect 211 341 269 347
rect 403 341 461 347
rect 595 341 653 347
rect 787 341 845 347
rect 979 341 1037 347
rect 1171 341 1229 347
rect 1363 341 1421 347
rect 1555 341 1613 347
rect 1747 341 1805 347
rect -1805 71 -1747 77
rect -1613 71 -1555 77
rect -1421 71 -1363 77
rect -1229 71 -1171 77
rect -1037 71 -979 77
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect 1075 71 1133 77
rect 1267 71 1325 77
rect 1459 71 1517 77
rect 1651 71 1709 77
rect 1843 71 1901 77
rect -1805 37 -1793 71
rect -1613 37 -1601 71
rect -1421 37 -1409 71
rect -1229 37 -1217 71
rect -1037 37 -1025 71
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect 1075 37 1087 71
rect 1267 37 1279 71
rect 1459 37 1471 71
rect 1651 37 1663 71
rect 1843 37 1855 71
rect -1805 31 -1747 37
rect -1613 31 -1555 37
rect -1421 31 -1363 37
rect -1229 31 -1171 37
rect -1037 31 -979 37
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect 1075 31 1133 37
rect 1267 31 1325 37
rect 1459 31 1517 37
rect 1651 31 1709 37
rect 1843 31 1901 37
rect -1805 -37 -1747 -31
rect -1613 -37 -1555 -31
rect -1421 -37 -1363 -31
rect -1229 -37 -1171 -31
rect -1037 -37 -979 -31
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect 1075 -37 1133 -31
rect 1267 -37 1325 -31
rect 1459 -37 1517 -31
rect 1651 -37 1709 -31
rect 1843 -37 1901 -31
rect -1805 -71 -1793 -37
rect -1613 -71 -1601 -37
rect -1421 -71 -1409 -37
rect -1229 -71 -1217 -37
rect -1037 -71 -1025 -37
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect 1075 -71 1087 -37
rect 1267 -71 1279 -37
rect 1459 -71 1471 -37
rect 1651 -71 1663 -37
rect 1843 -71 1855 -37
rect -1805 -77 -1747 -71
rect -1613 -77 -1555 -71
rect -1421 -77 -1363 -71
rect -1229 -77 -1171 -71
rect -1037 -77 -979 -71
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect 1075 -77 1133 -71
rect 1267 -77 1325 -71
rect 1459 -77 1517 -71
rect 1651 -77 1709 -71
rect 1843 -77 1901 -71
rect -1901 -347 -1843 -341
rect -1709 -347 -1651 -341
rect -1517 -347 -1459 -341
rect -1325 -347 -1267 -341
rect -1133 -347 -1075 -341
rect -941 -347 -883 -341
rect -749 -347 -691 -341
rect -557 -347 -499 -341
rect -365 -347 -307 -341
rect -173 -347 -115 -341
rect 19 -347 77 -341
rect 211 -347 269 -341
rect 403 -347 461 -341
rect 595 -347 653 -341
rect 787 -347 845 -341
rect 979 -347 1037 -341
rect 1171 -347 1229 -341
rect 1363 -347 1421 -341
rect 1555 -347 1613 -341
rect 1747 -347 1805 -341
rect -1901 -381 -1889 -347
rect -1709 -381 -1697 -347
rect -1517 -381 -1505 -347
rect -1325 -381 -1313 -347
rect -1133 -381 -1121 -347
rect -941 -381 -929 -347
rect -749 -381 -737 -347
rect -557 -381 -545 -347
rect -365 -381 -353 -347
rect -173 -381 -161 -347
rect 19 -381 31 -347
rect 211 -381 223 -347
rect 403 -381 415 -347
rect 595 -381 607 -347
rect 787 -381 799 -347
rect 979 -381 991 -347
rect 1171 -381 1183 -347
rect 1363 -381 1375 -347
rect 1555 -381 1567 -347
rect 1747 -381 1759 -347
rect -1901 -387 -1843 -381
rect -1709 -387 -1651 -381
rect -1517 -387 -1459 -381
rect -1325 -387 -1267 -381
rect -1133 -387 -1075 -381
rect -941 -387 -883 -381
rect -749 -387 -691 -381
rect -557 -387 -499 -381
rect -365 -387 -307 -381
rect -173 -387 -115 -381
rect 19 -387 77 -381
rect 211 -387 269 -381
rect 403 -387 461 -381
rect 595 -387 653 -381
rect 787 -387 845 -381
rect 979 -387 1037 -381
rect 1171 -387 1229 -381
rect 1363 -387 1421 -381
rect 1555 -387 1613 -381
rect 1747 -387 1805 -381
<< pwell >>
rect -2087 -519 2087 519
<< nmos >>
rect -1887 109 -1857 309
rect -1791 109 -1761 309
rect -1695 109 -1665 309
rect -1599 109 -1569 309
rect -1503 109 -1473 309
rect -1407 109 -1377 309
rect -1311 109 -1281 309
rect -1215 109 -1185 309
rect -1119 109 -1089 309
rect -1023 109 -993 309
rect -927 109 -897 309
rect -831 109 -801 309
rect -735 109 -705 309
rect -639 109 -609 309
rect -543 109 -513 309
rect -447 109 -417 309
rect -351 109 -321 309
rect -255 109 -225 309
rect -159 109 -129 309
rect -63 109 -33 309
rect 33 109 63 309
rect 129 109 159 309
rect 225 109 255 309
rect 321 109 351 309
rect 417 109 447 309
rect 513 109 543 309
rect 609 109 639 309
rect 705 109 735 309
rect 801 109 831 309
rect 897 109 927 309
rect 993 109 1023 309
rect 1089 109 1119 309
rect 1185 109 1215 309
rect 1281 109 1311 309
rect 1377 109 1407 309
rect 1473 109 1503 309
rect 1569 109 1599 309
rect 1665 109 1695 309
rect 1761 109 1791 309
rect 1857 109 1887 309
rect -1887 -309 -1857 -109
rect -1791 -309 -1761 -109
rect -1695 -309 -1665 -109
rect -1599 -309 -1569 -109
rect -1503 -309 -1473 -109
rect -1407 -309 -1377 -109
rect -1311 -309 -1281 -109
rect -1215 -309 -1185 -109
rect -1119 -309 -1089 -109
rect -1023 -309 -993 -109
rect -927 -309 -897 -109
rect -831 -309 -801 -109
rect -735 -309 -705 -109
rect -639 -309 -609 -109
rect -543 -309 -513 -109
rect -447 -309 -417 -109
rect -351 -309 -321 -109
rect -255 -309 -225 -109
rect -159 -309 -129 -109
rect -63 -309 -33 -109
rect 33 -309 63 -109
rect 129 -309 159 -109
rect 225 -309 255 -109
rect 321 -309 351 -109
rect 417 -309 447 -109
rect 513 -309 543 -109
rect 609 -309 639 -109
rect 705 -309 735 -109
rect 801 -309 831 -109
rect 897 -309 927 -109
rect 993 -309 1023 -109
rect 1089 -309 1119 -109
rect 1185 -309 1215 -109
rect 1281 -309 1311 -109
rect 1377 -309 1407 -109
rect 1473 -309 1503 -109
rect 1569 -309 1599 -109
rect 1665 -309 1695 -109
rect 1761 -309 1791 -109
rect 1857 -309 1887 -109
<< ndiff >>
rect -1949 297 -1887 309
rect -1949 121 -1937 297
rect -1903 121 -1887 297
rect -1949 109 -1887 121
rect -1857 297 -1791 309
rect -1857 121 -1841 297
rect -1807 121 -1791 297
rect -1857 109 -1791 121
rect -1761 297 -1695 309
rect -1761 121 -1745 297
rect -1711 121 -1695 297
rect -1761 109 -1695 121
rect -1665 297 -1599 309
rect -1665 121 -1649 297
rect -1615 121 -1599 297
rect -1665 109 -1599 121
rect -1569 297 -1503 309
rect -1569 121 -1553 297
rect -1519 121 -1503 297
rect -1569 109 -1503 121
rect -1473 297 -1407 309
rect -1473 121 -1457 297
rect -1423 121 -1407 297
rect -1473 109 -1407 121
rect -1377 297 -1311 309
rect -1377 121 -1361 297
rect -1327 121 -1311 297
rect -1377 109 -1311 121
rect -1281 297 -1215 309
rect -1281 121 -1265 297
rect -1231 121 -1215 297
rect -1281 109 -1215 121
rect -1185 297 -1119 309
rect -1185 121 -1169 297
rect -1135 121 -1119 297
rect -1185 109 -1119 121
rect -1089 297 -1023 309
rect -1089 121 -1073 297
rect -1039 121 -1023 297
rect -1089 109 -1023 121
rect -993 297 -927 309
rect -993 121 -977 297
rect -943 121 -927 297
rect -993 109 -927 121
rect -897 297 -831 309
rect -897 121 -881 297
rect -847 121 -831 297
rect -897 109 -831 121
rect -801 297 -735 309
rect -801 121 -785 297
rect -751 121 -735 297
rect -801 109 -735 121
rect -705 297 -639 309
rect -705 121 -689 297
rect -655 121 -639 297
rect -705 109 -639 121
rect -609 297 -543 309
rect -609 121 -593 297
rect -559 121 -543 297
rect -609 109 -543 121
rect -513 297 -447 309
rect -513 121 -497 297
rect -463 121 -447 297
rect -513 109 -447 121
rect -417 297 -351 309
rect -417 121 -401 297
rect -367 121 -351 297
rect -417 109 -351 121
rect -321 297 -255 309
rect -321 121 -305 297
rect -271 121 -255 297
rect -321 109 -255 121
rect -225 297 -159 309
rect -225 121 -209 297
rect -175 121 -159 297
rect -225 109 -159 121
rect -129 297 -63 309
rect -129 121 -113 297
rect -79 121 -63 297
rect -129 109 -63 121
rect -33 297 33 309
rect -33 121 -17 297
rect 17 121 33 297
rect -33 109 33 121
rect 63 297 129 309
rect 63 121 79 297
rect 113 121 129 297
rect 63 109 129 121
rect 159 297 225 309
rect 159 121 175 297
rect 209 121 225 297
rect 159 109 225 121
rect 255 297 321 309
rect 255 121 271 297
rect 305 121 321 297
rect 255 109 321 121
rect 351 297 417 309
rect 351 121 367 297
rect 401 121 417 297
rect 351 109 417 121
rect 447 297 513 309
rect 447 121 463 297
rect 497 121 513 297
rect 447 109 513 121
rect 543 297 609 309
rect 543 121 559 297
rect 593 121 609 297
rect 543 109 609 121
rect 639 297 705 309
rect 639 121 655 297
rect 689 121 705 297
rect 639 109 705 121
rect 735 297 801 309
rect 735 121 751 297
rect 785 121 801 297
rect 735 109 801 121
rect 831 297 897 309
rect 831 121 847 297
rect 881 121 897 297
rect 831 109 897 121
rect 927 297 993 309
rect 927 121 943 297
rect 977 121 993 297
rect 927 109 993 121
rect 1023 297 1089 309
rect 1023 121 1039 297
rect 1073 121 1089 297
rect 1023 109 1089 121
rect 1119 297 1185 309
rect 1119 121 1135 297
rect 1169 121 1185 297
rect 1119 109 1185 121
rect 1215 297 1281 309
rect 1215 121 1231 297
rect 1265 121 1281 297
rect 1215 109 1281 121
rect 1311 297 1377 309
rect 1311 121 1327 297
rect 1361 121 1377 297
rect 1311 109 1377 121
rect 1407 297 1473 309
rect 1407 121 1423 297
rect 1457 121 1473 297
rect 1407 109 1473 121
rect 1503 297 1569 309
rect 1503 121 1519 297
rect 1553 121 1569 297
rect 1503 109 1569 121
rect 1599 297 1665 309
rect 1599 121 1615 297
rect 1649 121 1665 297
rect 1599 109 1665 121
rect 1695 297 1761 309
rect 1695 121 1711 297
rect 1745 121 1761 297
rect 1695 109 1761 121
rect 1791 297 1857 309
rect 1791 121 1807 297
rect 1841 121 1857 297
rect 1791 109 1857 121
rect 1887 297 1949 309
rect 1887 121 1903 297
rect 1937 121 1949 297
rect 1887 109 1949 121
rect -1949 -121 -1887 -109
rect -1949 -297 -1937 -121
rect -1903 -297 -1887 -121
rect -1949 -309 -1887 -297
rect -1857 -121 -1791 -109
rect -1857 -297 -1841 -121
rect -1807 -297 -1791 -121
rect -1857 -309 -1791 -297
rect -1761 -121 -1695 -109
rect -1761 -297 -1745 -121
rect -1711 -297 -1695 -121
rect -1761 -309 -1695 -297
rect -1665 -121 -1599 -109
rect -1665 -297 -1649 -121
rect -1615 -297 -1599 -121
rect -1665 -309 -1599 -297
rect -1569 -121 -1503 -109
rect -1569 -297 -1553 -121
rect -1519 -297 -1503 -121
rect -1569 -309 -1503 -297
rect -1473 -121 -1407 -109
rect -1473 -297 -1457 -121
rect -1423 -297 -1407 -121
rect -1473 -309 -1407 -297
rect -1377 -121 -1311 -109
rect -1377 -297 -1361 -121
rect -1327 -297 -1311 -121
rect -1377 -309 -1311 -297
rect -1281 -121 -1215 -109
rect -1281 -297 -1265 -121
rect -1231 -297 -1215 -121
rect -1281 -309 -1215 -297
rect -1185 -121 -1119 -109
rect -1185 -297 -1169 -121
rect -1135 -297 -1119 -121
rect -1185 -309 -1119 -297
rect -1089 -121 -1023 -109
rect -1089 -297 -1073 -121
rect -1039 -297 -1023 -121
rect -1089 -309 -1023 -297
rect -993 -121 -927 -109
rect -993 -297 -977 -121
rect -943 -297 -927 -121
rect -993 -309 -927 -297
rect -897 -121 -831 -109
rect -897 -297 -881 -121
rect -847 -297 -831 -121
rect -897 -309 -831 -297
rect -801 -121 -735 -109
rect -801 -297 -785 -121
rect -751 -297 -735 -121
rect -801 -309 -735 -297
rect -705 -121 -639 -109
rect -705 -297 -689 -121
rect -655 -297 -639 -121
rect -705 -309 -639 -297
rect -609 -121 -543 -109
rect -609 -297 -593 -121
rect -559 -297 -543 -121
rect -609 -309 -543 -297
rect -513 -121 -447 -109
rect -513 -297 -497 -121
rect -463 -297 -447 -121
rect -513 -309 -447 -297
rect -417 -121 -351 -109
rect -417 -297 -401 -121
rect -367 -297 -351 -121
rect -417 -309 -351 -297
rect -321 -121 -255 -109
rect -321 -297 -305 -121
rect -271 -297 -255 -121
rect -321 -309 -255 -297
rect -225 -121 -159 -109
rect -225 -297 -209 -121
rect -175 -297 -159 -121
rect -225 -309 -159 -297
rect -129 -121 -63 -109
rect -129 -297 -113 -121
rect -79 -297 -63 -121
rect -129 -309 -63 -297
rect -33 -121 33 -109
rect -33 -297 -17 -121
rect 17 -297 33 -121
rect -33 -309 33 -297
rect 63 -121 129 -109
rect 63 -297 79 -121
rect 113 -297 129 -121
rect 63 -309 129 -297
rect 159 -121 225 -109
rect 159 -297 175 -121
rect 209 -297 225 -121
rect 159 -309 225 -297
rect 255 -121 321 -109
rect 255 -297 271 -121
rect 305 -297 321 -121
rect 255 -309 321 -297
rect 351 -121 417 -109
rect 351 -297 367 -121
rect 401 -297 417 -121
rect 351 -309 417 -297
rect 447 -121 513 -109
rect 447 -297 463 -121
rect 497 -297 513 -121
rect 447 -309 513 -297
rect 543 -121 609 -109
rect 543 -297 559 -121
rect 593 -297 609 -121
rect 543 -309 609 -297
rect 639 -121 705 -109
rect 639 -297 655 -121
rect 689 -297 705 -121
rect 639 -309 705 -297
rect 735 -121 801 -109
rect 735 -297 751 -121
rect 785 -297 801 -121
rect 735 -309 801 -297
rect 831 -121 897 -109
rect 831 -297 847 -121
rect 881 -297 897 -121
rect 831 -309 897 -297
rect 927 -121 993 -109
rect 927 -297 943 -121
rect 977 -297 993 -121
rect 927 -309 993 -297
rect 1023 -121 1089 -109
rect 1023 -297 1039 -121
rect 1073 -297 1089 -121
rect 1023 -309 1089 -297
rect 1119 -121 1185 -109
rect 1119 -297 1135 -121
rect 1169 -297 1185 -121
rect 1119 -309 1185 -297
rect 1215 -121 1281 -109
rect 1215 -297 1231 -121
rect 1265 -297 1281 -121
rect 1215 -309 1281 -297
rect 1311 -121 1377 -109
rect 1311 -297 1327 -121
rect 1361 -297 1377 -121
rect 1311 -309 1377 -297
rect 1407 -121 1473 -109
rect 1407 -297 1423 -121
rect 1457 -297 1473 -121
rect 1407 -309 1473 -297
rect 1503 -121 1569 -109
rect 1503 -297 1519 -121
rect 1553 -297 1569 -121
rect 1503 -309 1569 -297
rect 1599 -121 1665 -109
rect 1599 -297 1615 -121
rect 1649 -297 1665 -121
rect 1599 -309 1665 -297
rect 1695 -121 1761 -109
rect 1695 -297 1711 -121
rect 1745 -297 1761 -121
rect 1695 -309 1761 -297
rect 1791 -121 1857 -109
rect 1791 -297 1807 -121
rect 1841 -297 1857 -121
rect 1791 -309 1857 -297
rect 1887 -121 1949 -109
rect 1887 -297 1903 -121
rect 1937 -297 1949 -121
rect 1887 -309 1949 -297
<< ndiffc >>
rect -1937 121 -1903 297
rect -1841 121 -1807 297
rect -1745 121 -1711 297
rect -1649 121 -1615 297
rect -1553 121 -1519 297
rect -1457 121 -1423 297
rect -1361 121 -1327 297
rect -1265 121 -1231 297
rect -1169 121 -1135 297
rect -1073 121 -1039 297
rect -977 121 -943 297
rect -881 121 -847 297
rect -785 121 -751 297
rect -689 121 -655 297
rect -593 121 -559 297
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect 559 121 593 297
rect 655 121 689 297
rect 751 121 785 297
rect 847 121 881 297
rect 943 121 977 297
rect 1039 121 1073 297
rect 1135 121 1169 297
rect 1231 121 1265 297
rect 1327 121 1361 297
rect 1423 121 1457 297
rect 1519 121 1553 297
rect 1615 121 1649 297
rect 1711 121 1745 297
rect 1807 121 1841 297
rect 1903 121 1937 297
rect -1937 -297 -1903 -121
rect -1841 -297 -1807 -121
rect -1745 -297 -1711 -121
rect -1649 -297 -1615 -121
rect -1553 -297 -1519 -121
rect -1457 -297 -1423 -121
rect -1361 -297 -1327 -121
rect -1265 -297 -1231 -121
rect -1169 -297 -1135 -121
rect -1073 -297 -1039 -121
rect -977 -297 -943 -121
rect -881 -297 -847 -121
rect -785 -297 -751 -121
rect -689 -297 -655 -121
rect -593 -297 -559 -121
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect 559 -297 593 -121
rect 655 -297 689 -121
rect 751 -297 785 -121
rect 847 -297 881 -121
rect 943 -297 977 -121
rect 1039 -297 1073 -121
rect 1135 -297 1169 -121
rect 1231 -297 1265 -121
rect 1327 -297 1361 -121
rect 1423 -297 1457 -121
rect 1519 -297 1553 -121
rect 1615 -297 1649 -121
rect 1711 -297 1745 -121
rect 1807 -297 1841 -121
rect 1903 -297 1937 -121
<< psubdiff >>
rect -2051 449 -1955 483
rect 1955 449 2051 483
rect -2051 387 -2017 449
rect 2017 387 2051 449
rect -2051 -449 -2017 -387
rect 2017 -449 2051 -387
rect -2051 -483 -1955 -449
rect 1955 -483 2051 -449
<< psubdiffcont >>
rect -1955 449 1955 483
rect -2051 -387 -2017 387
rect 2017 -387 2051 387
rect -1955 -483 1955 -449
<< poly >>
rect -1905 381 -1839 397
rect -1905 347 -1889 381
rect -1855 347 -1839 381
rect -1905 331 -1839 347
rect -1713 381 -1647 397
rect -1713 347 -1697 381
rect -1663 347 -1647 381
rect -1887 309 -1857 331
rect -1791 309 -1761 335
rect -1713 331 -1647 347
rect -1521 381 -1455 397
rect -1521 347 -1505 381
rect -1471 347 -1455 381
rect -1695 309 -1665 331
rect -1599 309 -1569 335
rect -1521 331 -1455 347
rect -1329 381 -1263 397
rect -1329 347 -1313 381
rect -1279 347 -1263 381
rect -1503 309 -1473 331
rect -1407 309 -1377 335
rect -1329 331 -1263 347
rect -1137 381 -1071 397
rect -1137 347 -1121 381
rect -1087 347 -1071 381
rect -1311 309 -1281 331
rect -1215 309 -1185 335
rect -1137 331 -1071 347
rect -945 381 -879 397
rect -945 347 -929 381
rect -895 347 -879 381
rect -1119 309 -1089 331
rect -1023 309 -993 335
rect -945 331 -879 347
rect -753 381 -687 397
rect -753 347 -737 381
rect -703 347 -687 381
rect -927 309 -897 331
rect -831 309 -801 335
rect -753 331 -687 347
rect -561 381 -495 397
rect -561 347 -545 381
rect -511 347 -495 381
rect -735 309 -705 331
rect -639 309 -609 335
rect -561 331 -495 347
rect -369 381 -303 397
rect -369 347 -353 381
rect -319 347 -303 381
rect -543 309 -513 331
rect -447 309 -417 335
rect -369 331 -303 347
rect -177 381 -111 397
rect -177 347 -161 381
rect -127 347 -111 381
rect -351 309 -321 331
rect -255 309 -225 335
rect -177 331 -111 347
rect 15 381 81 397
rect 15 347 31 381
rect 65 347 81 381
rect -159 309 -129 331
rect -63 309 -33 335
rect 15 331 81 347
rect 207 381 273 397
rect 207 347 223 381
rect 257 347 273 381
rect 33 309 63 331
rect 129 309 159 335
rect 207 331 273 347
rect 399 381 465 397
rect 399 347 415 381
rect 449 347 465 381
rect 225 309 255 331
rect 321 309 351 335
rect 399 331 465 347
rect 591 381 657 397
rect 591 347 607 381
rect 641 347 657 381
rect 417 309 447 331
rect 513 309 543 335
rect 591 331 657 347
rect 783 381 849 397
rect 783 347 799 381
rect 833 347 849 381
rect 609 309 639 331
rect 705 309 735 335
rect 783 331 849 347
rect 975 381 1041 397
rect 975 347 991 381
rect 1025 347 1041 381
rect 801 309 831 331
rect 897 309 927 335
rect 975 331 1041 347
rect 1167 381 1233 397
rect 1167 347 1183 381
rect 1217 347 1233 381
rect 993 309 1023 331
rect 1089 309 1119 335
rect 1167 331 1233 347
rect 1359 381 1425 397
rect 1359 347 1375 381
rect 1409 347 1425 381
rect 1185 309 1215 331
rect 1281 309 1311 335
rect 1359 331 1425 347
rect 1551 381 1617 397
rect 1551 347 1567 381
rect 1601 347 1617 381
rect 1377 309 1407 331
rect 1473 309 1503 335
rect 1551 331 1617 347
rect 1743 381 1809 397
rect 1743 347 1759 381
rect 1793 347 1809 381
rect 1569 309 1599 331
rect 1665 309 1695 335
rect 1743 331 1809 347
rect 1761 309 1791 331
rect 1857 309 1887 335
rect -1887 83 -1857 109
rect -1791 87 -1761 109
rect -1809 71 -1743 87
rect -1695 83 -1665 109
rect -1599 87 -1569 109
rect -1809 37 -1793 71
rect -1759 37 -1743 71
rect -1809 21 -1743 37
rect -1617 71 -1551 87
rect -1503 83 -1473 109
rect -1407 87 -1377 109
rect -1617 37 -1601 71
rect -1567 37 -1551 71
rect -1617 21 -1551 37
rect -1425 71 -1359 87
rect -1311 83 -1281 109
rect -1215 87 -1185 109
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1425 21 -1359 37
rect -1233 71 -1167 87
rect -1119 83 -1089 109
rect -1023 87 -993 109
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1233 21 -1167 37
rect -1041 71 -975 87
rect -927 83 -897 109
rect -831 87 -801 109
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -1041 21 -975 37
rect -849 71 -783 87
rect -735 83 -705 109
rect -639 87 -609 109
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -543 83 -513 109
rect -447 87 -417 109
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -351 83 -321 109
rect -255 87 -225 109
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -159 83 -129 109
rect -63 87 -33 109
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 225 83 255 109
rect 321 87 351 109
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 417 83 447 109
rect 513 87 543 109
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 609 83 639 109
rect 705 87 735 109
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 801 83 831 109
rect 897 87 927 109
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 993 83 1023 109
rect 1089 87 1119 109
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect 1071 71 1137 87
rect 1185 83 1215 109
rect 1281 87 1311 109
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1071 21 1137 37
rect 1263 71 1329 87
rect 1377 83 1407 109
rect 1473 87 1503 109
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1263 21 1329 37
rect 1455 71 1521 87
rect 1569 83 1599 109
rect 1665 87 1695 109
rect 1455 37 1471 71
rect 1505 37 1521 71
rect 1455 21 1521 37
rect 1647 71 1713 87
rect 1761 83 1791 109
rect 1857 87 1887 109
rect 1647 37 1663 71
rect 1697 37 1713 71
rect 1647 21 1713 37
rect 1839 71 1905 87
rect 1839 37 1855 71
rect 1889 37 1905 71
rect 1839 21 1905 37
rect -1809 -37 -1743 -21
rect -1809 -71 -1793 -37
rect -1759 -71 -1743 -37
rect -1887 -109 -1857 -83
rect -1809 -87 -1743 -71
rect -1617 -37 -1551 -21
rect -1617 -71 -1601 -37
rect -1567 -71 -1551 -37
rect -1791 -109 -1761 -87
rect -1695 -109 -1665 -83
rect -1617 -87 -1551 -71
rect -1425 -37 -1359 -21
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1599 -109 -1569 -87
rect -1503 -109 -1473 -83
rect -1425 -87 -1359 -71
rect -1233 -37 -1167 -21
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1407 -109 -1377 -87
rect -1311 -109 -1281 -83
rect -1233 -87 -1167 -71
rect -1041 -37 -975 -21
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -1215 -109 -1185 -87
rect -1119 -109 -1089 -83
rect -1041 -87 -975 -71
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -1023 -109 -993 -87
rect -927 -109 -897 -83
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -831 -109 -801 -87
rect -735 -109 -705 -83
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -639 -109 -609 -87
rect -543 -109 -513 -83
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -447 -109 -417 -87
rect -351 -109 -321 -83
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -255 -109 -225 -87
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 129 -109 159 -87
rect 225 -109 255 -83
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 321 -109 351 -87
rect 417 -109 447 -83
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 513 -109 543 -87
rect 609 -109 639 -83
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 705 -109 735 -87
rect 801 -109 831 -83
rect 879 -87 945 -71
rect 1071 -37 1137 -21
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 897 -109 927 -87
rect 993 -109 1023 -83
rect 1071 -87 1137 -71
rect 1263 -37 1329 -21
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1089 -109 1119 -87
rect 1185 -109 1215 -83
rect 1263 -87 1329 -71
rect 1455 -37 1521 -21
rect 1455 -71 1471 -37
rect 1505 -71 1521 -37
rect 1281 -109 1311 -87
rect 1377 -109 1407 -83
rect 1455 -87 1521 -71
rect 1647 -37 1713 -21
rect 1647 -71 1663 -37
rect 1697 -71 1713 -37
rect 1473 -109 1503 -87
rect 1569 -109 1599 -83
rect 1647 -87 1713 -71
rect 1839 -37 1905 -21
rect 1839 -71 1855 -37
rect 1889 -71 1905 -37
rect 1665 -109 1695 -87
rect 1761 -109 1791 -83
rect 1839 -87 1905 -71
rect 1857 -109 1887 -87
rect -1887 -331 -1857 -309
rect -1905 -347 -1839 -331
rect -1791 -335 -1761 -309
rect -1695 -331 -1665 -309
rect -1905 -381 -1889 -347
rect -1855 -381 -1839 -347
rect -1905 -397 -1839 -381
rect -1713 -347 -1647 -331
rect -1599 -335 -1569 -309
rect -1503 -331 -1473 -309
rect -1713 -381 -1697 -347
rect -1663 -381 -1647 -347
rect -1713 -397 -1647 -381
rect -1521 -347 -1455 -331
rect -1407 -335 -1377 -309
rect -1311 -331 -1281 -309
rect -1521 -381 -1505 -347
rect -1471 -381 -1455 -347
rect -1521 -397 -1455 -381
rect -1329 -347 -1263 -331
rect -1215 -335 -1185 -309
rect -1119 -331 -1089 -309
rect -1329 -381 -1313 -347
rect -1279 -381 -1263 -347
rect -1329 -397 -1263 -381
rect -1137 -347 -1071 -331
rect -1023 -335 -993 -309
rect -927 -331 -897 -309
rect -1137 -381 -1121 -347
rect -1087 -381 -1071 -347
rect -1137 -397 -1071 -381
rect -945 -347 -879 -331
rect -831 -335 -801 -309
rect -735 -331 -705 -309
rect -945 -381 -929 -347
rect -895 -381 -879 -347
rect -945 -397 -879 -381
rect -753 -347 -687 -331
rect -639 -335 -609 -309
rect -543 -331 -513 -309
rect -753 -381 -737 -347
rect -703 -381 -687 -347
rect -753 -397 -687 -381
rect -561 -347 -495 -331
rect -447 -335 -417 -309
rect -351 -331 -321 -309
rect -561 -381 -545 -347
rect -511 -381 -495 -347
rect -561 -397 -495 -381
rect -369 -347 -303 -331
rect -255 -335 -225 -309
rect -159 -331 -129 -309
rect -369 -381 -353 -347
rect -319 -381 -303 -347
rect -369 -397 -303 -381
rect -177 -347 -111 -331
rect -63 -335 -33 -309
rect 33 -331 63 -309
rect -177 -381 -161 -347
rect -127 -381 -111 -347
rect -177 -397 -111 -381
rect 15 -347 81 -331
rect 129 -335 159 -309
rect 225 -331 255 -309
rect 15 -381 31 -347
rect 65 -381 81 -347
rect 15 -397 81 -381
rect 207 -347 273 -331
rect 321 -335 351 -309
rect 417 -331 447 -309
rect 207 -381 223 -347
rect 257 -381 273 -347
rect 207 -397 273 -381
rect 399 -347 465 -331
rect 513 -335 543 -309
rect 609 -331 639 -309
rect 399 -381 415 -347
rect 449 -381 465 -347
rect 399 -397 465 -381
rect 591 -347 657 -331
rect 705 -335 735 -309
rect 801 -331 831 -309
rect 591 -381 607 -347
rect 641 -381 657 -347
rect 591 -397 657 -381
rect 783 -347 849 -331
rect 897 -335 927 -309
rect 993 -331 1023 -309
rect 783 -381 799 -347
rect 833 -381 849 -347
rect 783 -397 849 -381
rect 975 -347 1041 -331
rect 1089 -335 1119 -309
rect 1185 -331 1215 -309
rect 975 -381 991 -347
rect 1025 -381 1041 -347
rect 975 -397 1041 -381
rect 1167 -347 1233 -331
rect 1281 -335 1311 -309
rect 1377 -331 1407 -309
rect 1167 -381 1183 -347
rect 1217 -381 1233 -347
rect 1167 -397 1233 -381
rect 1359 -347 1425 -331
rect 1473 -335 1503 -309
rect 1569 -331 1599 -309
rect 1359 -381 1375 -347
rect 1409 -381 1425 -347
rect 1359 -397 1425 -381
rect 1551 -347 1617 -331
rect 1665 -335 1695 -309
rect 1761 -331 1791 -309
rect 1551 -381 1567 -347
rect 1601 -381 1617 -347
rect 1551 -397 1617 -381
rect 1743 -347 1809 -331
rect 1857 -335 1887 -309
rect 1743 -381 1759 -347
rect 1793 -381 1809 -347
rect 1743 -397 1809 -381
<< polycont >>
rect -1889 347 -1855 381
rect -1697 347 -1663 381
rect -1505 347 -1471 381
rect -1313 347 -1279 381
rect -1121 347 -1087 381
rect -929 347 -895 381
rect -737 347 -703 381
rect -545 347 -511 381
rect -353 347 -319 381
rect -161 347 -127 381
rect 31 347 65 381
rect 223 347 257 381
rect 415 347 449 381
rect 607 347 641 381
rect 799 347 833 381
rect 991 347 1025 381
rect 1183 347 1217 381
rect 1375 347 1409 381
rect 1567 347 1601 381
rect 1759 347 1793 381
rect -1793 37 -1759 71
rect -1601 37 -1567 71
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect 1471 37 1505 71
rect 1663 37 1697 71
rect 1855 37 1889 71
rect -1793 -71 -1759 -37
rect -1601 -71 -1567 -37
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect 1471 -71 1505 -37
rect 1663 -71 1697 -37
rect 1855 -71 1889 -37
rect -1889 -381 -1855 -347
rect -1697 -381 -1663 -347
rect -1505 -381 -1471 -347
rect -1313 -381 -1279 -347
rect -1121 -381 -1087 -347
rect -929 -381 -895 -347
rect -737 -381 -703 -347
rect -545 -381 -511 -347
rect -353 -381 -319 -347
rect -161 -381 -127 -347
rect 31 -381 65 -347
rect 223 -381 257 -347
rect 415 -381 449 -347
rect 607 -381 641 -347
rect 799 -381 833 -347
rect 991 -381 1025 -347
rect 1183 -381 1217 -347
rect 1375 -381 1409 -347
rect 1567 -381 1601 -347
rect 1759 -381 1793 -347
<< locali >>
rect -2051 449 -1955 483
rect 1955 449 2051 483
rect -2051 387 -2017 449
rect 2017 387 2051 449
rect -1905 347 -1889 381
rect -1855 347 -1839 381
rect -1713 347 -1697 381
rect -1663 347 -1647 381
rect -1521 347 -1505 381
rect -1471 347 -1455 381
rect -1329 347 -1313 381
rect -1279 347 -1263 381
rect -1137 347 -1121 381
rect -1087 347 -1071 381
rect -945 347 -929 381
rect -895 347 -879 381
rect -753 347 -737 381
rect -703 347 -687 381
rect -561 347 -545 381
rect -511 347 -495 381
rect -369 347 -353 381
rect -319 347 -303 381
rect -177 347 -161 381
rect -127 347 -111 381
rect 15 347 31 381
rect 65 347 81 381
rect 207 347 223 381
rect 257 347 273 381
rect 399 347 415 381
rect 449 347 465 381
rect 591 347 607 381
rect 641 347 657 381
rect 783 347 799 381
rect 833 347 849 381
rect 975 347 991 381
rect 1025 347 1041 381
rect 1167 347 1183 381
rect 1217 347 1233 381
rect 1359 347 1375 381
rect 1409 347 1425 381
rect 1551 347 1567 381
rect 1601 347 1617 381
rect 1743 347 1759 381
rect 1793 347 1809 381
rect -1937 297 -1903 313
rect -1937 105 -1903 121
rect -1841 297 -1807 313
rect -1841 105 -1807 121
rect -1745 297 -1711 313
rect -1745 105 -1711 121
rect -1649 297 -1615 313
rect -1649 105 -1615 121
rect -1553 297 -1519 313
rect -1553 105 -1519 121
rect -1457 297 -1423 313
rect -1457 105 -1423 121
rect -1361 297 -1327 313
rect -1361 105 -1327 121
rect -1265 297 -1231 313
rect -1265 105 -1231 121
rect -1169 297 -1135 313
rect -1169 105 -1135 121
rect -1073 297 -1039 313
rect -1073 105 -1039 121
rect -977 297 -943 313
rect -977 105 -943 121
rect -881 297 -847 313
rect -881 105 -847 121
rect -785 297 -751 313
rect -785 105 -751 121
rect -689 297 -655 313
rect -689 105 -655 121
rect -593 297 -559 313
rect -593 105 -559 121
rect -497 297 -463 313
rect -497 105 -463 121
rect -401 297 -367 313
rect -401 105 -367 121
rect -305 297 -271 313
rect -305 105 -271 121
rect -209 297 -175 313
rect -209 105 -175 121
rect -113 297 -79 313
rect -113 105 -79 121
rect -17 297 17 313
rect -17 105 17 121
rect 79 297 113 313
rect 79 105 113 121
rect 175 297 209 313
rect 175 105 209 121
rect 271 297 305 313
rect 271 105 305 121
rect 367 297 401 313
rect 367 105 401 121
rect 463 297 497 313
rect 463 105 497 121
rect 559 297 593 313
rect 559 105 593 121
rect 655 297 689 313
rect 655 105 689 121
rect 751 297 785 313
rect 751 105 785 121
rect 847 297 881 313
rect 847 105 881 121
rect 943 297 977 313
rect 943 105 977 121
rect 1039 297 1073 313
rect 1039 105 1073 121
rect 1135 297 1169 313
rect 1135 105 1169 121
rect 1231 297 1265 313
rect 1231 105 1265 121
rect 1327 297 1361 313
rect 1327 105 1361 121
rect 1423 297 1457 313
rect 1423 105 1457 121
rect 1519 297 1553 313
rect 1519 105 1553 121
rect 1615 297 1649 313
rect 1615 105 1649 121
rect 1711 297 1745 313
rect 1711 105 1745 121
rect 1807 297 1841 313
rect 1807 105 1841 121
rect 1903 297 1937 313
rect 1903 105 1937 121
rect -1809 37 -1793 71
rect -1759 37 -1743 71
rect -1617 37 -1601 71
rect -1567 37 -1551 71
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1455 37 1471 71
rect 1505 37 1521 71
rect 1647 37 1663 71
rect 1697 37 1713 71
rect 1839 37 1855 71
rect 1889 37 1905 71
rect -1809 -71 -1793 -37
rect -1759 -71 -1743 -37
rect -1617 -71 -1601 -37
rect -1567 -71 -1551 -37
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1455 -71 1471 -37
rect 1505 -71 1521 -37
rect 1647 -71 1663 -37
rect 1697 -71 1713 -37
rect 1839 -71 1855 -37
rect 1889 -71 1905 -37
rect -1937 -121 -1903 -105
rect -1937 -313 -1903 -297
rect -1841 -121 -1807 -105
rect -1841 -313 -1807 -297
rect -1745 -121 -1711 -105
rect -1745 -313 -1711 -297
rect -1649 -121 -1615 -105
rect -1649 -313 -1615 -297
rect -1553 -121 -1519 -105
rect -1553 -313 -1519 -297
rect -1457 -121 -1423 -105
rect -1457 -313 -1423 -297
rect -1361 -121 -1327 -105
rect -1361 -313 -1327 -297
rect -1265 -121 -1231 -105
rect -1265 -313 -1231 -297
rect -1169 -121 -1135 -105
rect -1169 -313 -1135 -297
rect -1073 -121 -1039 -105
rect -1073 -313 -1039 -297
rect -977 -121 -943 -105
rect -977 -313 -943 -297
rect -881 -121 -847 -105
rect -881 -313 -847 -297
rect -785 -121 -751 -105
rect -785 -313 -751 -297
rect -689 -121 -655 -105
rect -689 -313 -655 -297
rect -593 -121 -559 -105
rect -593 -313 -559 -297
rect -497 -121 -463 -105
rect -497 -313 -463 -297
rect -401 -121 -367 -105
rect -401 -313 -367 -297
rect -305 -121 -271 -105
rect -305 -313 -271 -297
rect -209 -121 -175 -105
rect -209 -313 -175 -297
rect -113 -121 -79 -105
rect -113 -313 -79 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 79 -121 113 -105
rect 79 -313 113 -297
rect 175 -121 209 -105
rect 175 -313 209 -297
rect 271 -121 305 -105
rect 271 -313 305 -297
rect 367 -121 401 -105
rect 367 -313 401 -297
rect 463 -121 497 -105
rect 463 -313 497 -297
rect 559 -121 593 -105
rect 559 -313 593 -297
rect 655 -121 689 -105
rect 655 -313 689 -297
rect 751 -121 785 -105
rect 751 -313 785 -297
rect 847 -121 881 -105
rect 847 -313 881 -297
rect 943 -121 977 -105
rect 943 -313 977 -297
rect 1039 -121 1073 -105
rect 1039 -313 1073 -297
rect 1135 -121 1169 -105
rect 1135 -313 1169 -297
rect 1231 -121 1265 -105
rect 1231 -313 1265 -297
rect 1327 -121 1361 -105
rect 1327 -313 1361 -297
rect 1423 -121 1457 -105
rect 1423 -313 1457 -297
rect 1519 -121 1553 -105
rect 1519 -313 1553 -297
rect 1615 -121 1649 -105
rect 1615 -313 1649 -297
rect 1711 -121 1745 -105
rect 1711 -313 1745 -297
rect 1807 -121 1841 -105
rect 1807 -313 1841 -297
rect 1903 -121 1937 -105
rect 1903 -313 1937 -297
rect -1905 -381 -1889 -347
rect -1855 -381 -1839 -347
rect -1713 -381 -1697 -347
rect -1663 -381 -1647 -347
rect -1521 -381 -1505 -347
rect -1471 -381 -1455 -347
rect -1329 -381 -1313 -347
rect -1279 -381 -1263 -347
rect -1137 -381 -1121 -347
rect -1087 -381 -1071 -347
rect -945 -381 -929 -347
rect -895 -381 -879 -347
rect -753 -381 -737 -347
rect -703 -381 -687 -347
rect -561 -381 -545 -347
rect -511 -381 -495 -347
rect -369 -381 -353 -347
rect -319 -381 -303 -347
rect -177 -381 -161 -347
rect -127 -381 -111 -347
rect 15 -381 31 -347
rect 65 -381 81 -347
rect 207 -381 223 -347
rect 257 -381 273 -347
rect 399 -381 415 -347
rect 449 -381 465 -347
rect 591 -381 607 -347
rect 641 -381 657 -347
rect 783 -381 799 -347
rect 833 -381 849 -347
rect 975 -381 991 -347
rect 1025 -381 1041 -347
rect 1167 -381 1183 -347
rect 1217 -381 1233 -347
rect 1359 -381 1375 -347
rect 1409 -381 1425 -347
rect 1551 -381 1567 -347
rect 1601 -381 1617 -347
rect 1743 -381 1759 -347
rect 1793 -381 1809 -347
rect -2051 -449 -2017 -387
rect 2017 -449 2051 -387
rect -2051 -483 -1955 -449
rect 1955 -483 2051 -449
<< viali >>
rect -1889 347 -1855 381
rect -1697 347 -1663 381
rect -1505 347 -1471 381
rect -1313 347 -1279 381
rect -1121 347 -1087 381
rect -929 347 -895 381
rect -737 347 -703 381
rect -545 347 -511 381
rect -353 347 -319 381
rect -161 347 -127 381
rect 31 347 65 381
rect 223 347 257 381
rect 415 347 449 381
rect 607 347 641 381
rect 799 347 833 381
rect 991 347 1025 381
rect 1183 347 1217 381
rect 1375 347 1409 381
rect 1567 347 1601 381
rect 1759 347 1793 381
rect -1937 121 -1903 297
rect -1841 121 -1807 297
rect -1745 121 -1711 297
rect -1649 121 -1615 297
rect -1553 121 -1519 297
rect -1457 121 -1423 297
rect -1361 121 -1327 297
rect -1265 121 -1231 297
rect -1169 121 -1135 297
rect -1073 121 -1039 297
rect -977 121 -943 297
rect -881 121 -847 297
rect -785 121 -751 297
rect -689 121 -655 297
rect -593 121 -559 297
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect 559 121 593 297
rect 655 121 689 297
rect 751 121 785 297
rect 847 121 881 297
rect 943 121 977 297
rect 1039 121 1073 297
rect 1135 121 1169 297
rect 1231 121 1265 297
rect 1327 121 1361 297
rect 1423 121 1457 297
rect 1519 121 1553 297
rect 1615 121 1649 297
rect 1711 121 1745 297
rect 1807 121 1841 297
rect 1903 121 1937 297
rect -1793 37 -1759 71
rect -1601 37 -1567 71
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect 1471 37 1505 71
rect 1663 37 1697 71
rect 1855 37 1889 71
rect -1793 -71 -1759 -37
rect -1601 -71 -1567 -37
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect 1471 -71 1505 -37
rect 1663 -71 1697 -37
rect 1855 -71 1889 -37
rect -1937 -297 -1903 -121
rect -1841 -297 -1807 -121
rect -1745 -297 -1711 -121
rect -1649 -297 -1615 -121
rect -1553 -297 -1519 -121
rect -1457 -297 -1423 -121
rect -1361 -297 -1327 -121
rect -1265 -297 -1231 -121
rect -1169 -297 -1135 -121
rect -1073 -297 -1039 -121
rect -977 -297 -943 -121
rect -881 -297 -847 -121
rect -785 -297 -751 -121
rect -689 -297 -655 -121
rect -593 -297 -559 -121
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect 559 -297 593 -121
rect 655 -297 689 -121
rect 751 -297 785 -121
rect 847 -297 881 -121
rect 943 -297 977 -121
rect 1039 -297 1073 -121
rect 1135 -297 1169 -121
rect 1231 -297 1265 -121
rect 1327 -297 1361 -121
rect 1423 -297 1457 -121
rect 1519 -297 1553 -121
rect 1615 -297 1649 -121
rect 1711 -297 1745 -121
rect 1807 -297 1841 -121
rect 1903 -297 1937 -121
rect -1889 -381 -1855 -347
rect -1697 -381 -1663 -347
rect -1505 -381 -1471 -347
rect -1313 -381 -1279 -347
rect -1121 -381 -1087 -347
rect -929 -381 -895 -347
rect -737 -381 -703 -347
rect -545 -381 -511 -347
rect -353 -381 -319 -347
rect -161 -381 -127 -347
rect 31 -381 65 -347
rect 223 -381 257 -347
rect 415 -381 449 -347
rect 607 -381 641 -347
rect 799 -381 833 -347
rect 991 -381 1025 -347
rect 1183 -381 1217 -347
rect 1375 -381 1409 -347
rect 1567 -381 1601 -347
rect 1759 -381 1793 -347
<< metal1 >>
rect -1901 381 -1843 387
rect -1901 347 -1889 381
rect -1855 347 -1843 381
rect -1901 341 -1843 347
rect -1709 381 -1651 387
rect -1709 347 -1697 381
rect -1663 347 -1651 381
rect -1709 341 -1651 347
rect -1517 381 -1459 387
rect -1517 347 -1505 381
rect -1471 347 -1459 381
rect -1517 341 -1459 347
rect -1325 381 -1267 387
rect -1325 347 -1313 381
rect -1279 347 -1267 381
rect -1325 341 -1267 347
rect -1133 381 -1075 387
rect -1133 347 -1121 381
rect -1087 347 -1075 381
rect -1133 341 -1075 347
rect -941 381 -883 387
rect -941 347 -929 381
rect -895 347 -883 381
rect -941 341 -883 347
rect -749 381 -691 387
rect -749 347 -737 381
rect -703 347 -691 381
rect -749 341 -691 347
rect -557 381 -499 387
rect -557 347 -545 381
rect -511 347 -499 381
rect -557 341 -499 347
rect -365 381 -307 387
rect -365 347 -353 381
rect -319 347 -307 381
rect -365 341 -307 347
rect -173 381 -115 387
rect -173 347 -161 381
rect -127 347 -115 381
rect -173 341 -115 347
rect 19 381 77 387
rect 19 347 31 381
rect 65 347 77 381
rect 19 341 77 347
rect 211 381 269 387
rect 211 347 223 381
rect 257 347 269 381
rect 211 341 269 347
rect 403 381 461 387
rect 403 347 415 381
rect 449 347 461 381
rect 403 341 461 347
rect 595 381 653 387
rect 595 347 607 381
rect 641 347 653 381
rect 595 341 653 347
rect 787 381 845 387
rect 787 347 799 381
rect 833 347 845 381
rect 787 341 845 347
rect 979 381 1037 387
rect 979 347 991 381
rect 1025 347 1037 381
rect 979 341 1037 347
rect 1171 381 1229 387
rect 1171 347 1183 381
rect 1217 347 1229 381
rect 1171 341 1229 347
rect 1363 381 1421 387
rect 1363 347 1375 381
rect 1409 347 1421 381
rect 1363 341 1421 347
rect 1555 381 1613 387
rect 1555 347 1567 381
rect 1601 347 1613 381
rect 1555 341 1613 347
rect 1747 381 1805 387
rect 1747 347 1759 381
rect 1793 347 1805 381
rect 1747 341 1805 347
rect -1943 297 -1897 309
rect -1943 121 -1937 297
rect -1903 121 -1897 297
rect -1943 109 -1897 121
rect -1847 297 -1801 309
rect -1847 121 -1841 297
rect -1807 121 -1801 297
rect -1847 109 -1801 121
rect -1751 297 -1705 309
rect -1751 121 -1745 297
rect -1711 121 -1705 297
rect -1751 109 -1705 121
rect -1655 297 -1609 309
rect -1655 121 -1649 297
rect -1615 121 -1609 297
rect -1655 109 -1609 121
rect -1559 297 -1513 309
rect -1559 121 -1553 297
rect -1519 121 -1513 297
rect -1559 109 -1513 121
rect -1463 297 -1417 309
rect -1463 121 -1457 297
rect -1423 121 -1417 297
rect -1463 109 -1417 121
rect -1367 297 -1321 309
rect -1367 121 -1361 297
rect -1327 121 -1321 297
rect -1367 109 -1321 121
rect -1271 297 -1225 309
rect -1271 121 -1265 297
rect -1231 121 -1225 297
rect -1271 109 -1225 121
rect -1175 297 -1129 309
rect -1175 121 -1169 297
rect -1135 121 -1129 297
rect -1175 109 -1129 121
rect -1079 297 -1033 309
rect -1079 121 -1073 297
rect -1039 121 -1033 297
rect -1079 109 -1033 121
rect -983 297 -937 309
rect -983 121 -977 297
rect -943 121 -937 297
rect -983 109 -937 121
rect -887 297 -841 309
rect -887 121 -881 297
rect -847 121 -841 297
rect -887 109 -841 121
rect -791 297 -745 309
rect -791 121 -785 297
rect -751 121 -745 297
rect -791 109 -745 121
rect -695 297 -649 309
rect -695 121 -689 297
rect -655 121 -649 297
rect -695 109 -649 121
rect -599 297 -553 309
rect -599 121 -593 297
rect -559 121 -553 297
rect -599 109 -553 121
rect -503 297 -457 309
rect -503 121 -497 297
rect -463 121 -457 297
rect -503 109 -457 121
rect -407 297 -361 309
rect -407 121 -401 297
rect -367 121 -361 297
rect -407 109 -361 121
rect -311 297 -265 309
rect -311 121 -305 297
rect -271 121 -265 297
rect -311 109 -265 121
rect -215 297 -169 309
rect -215 121 -209 297
rect -175 121 -169 297
rect -215 109 -169 121
rect -119 297 -73 309
rect -119 121 -113 297
rect -79 121 -73 297
rect -119 109 -73 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 73 297 119 309
rect 73 121 79 297
rect 113 121 119 297
rect 73 109 119 121
rect 169 297 215 309
rect 169 121 175 297
rect 209 121 215 297
rect 169 109 215 121
rect 265 297 311 309
rect 265 121 271 297
rect 305 121 311 297
rect 265 109 311 121
rect 361 297 407 309
rect 361 121 367 297
rect 401 121 407 297
rect 361 109 407 121
rect 457 297 503 309
rect 457 121 463 297
rect 497 121 503 297
rect 457 109 503 121
rect 553 297 599 309
rect 553 121 559 297
rect 593 121 599 297
rect 553 109 599 121
rect 649 297 695 309
rect 649 121 655 297
rect 689 121 695 297
rect 649 109 695 121
rect 745 297 791 309
rect 745 121 751 297
rect 785 121 791 297
rect 745 109 791 121
rect 841 297 887 309
rect 841 121 847 297
rect 881 121 887 297
rect 841 109 887 121
rect 937 297 983 309
rect 937 121 943 297
rect 977 121 983 297
rect 937 109 983 121
rect 1033 297 1079 309
rect 1033 121 1039 297
rect 1073 121 1079 297
rect 1033 109 1079 121
rect 1129 297 1175 309
rect 1129 121 1135 297
rect 1169 121 1175 297
rect 1129 109 1175 121
rect 1225 297 1271 309
rect 1225 121 1231 297
rect 1265 121 1271 297
rect 1225 109 1271 121
rect 1321 297 1367 309
rect 1321 121 1327 297
rect 1361 121 1367 297
rect 1321 109 1367 121
rect 1417 297 1463 309
rect 1417 121 1423 297
rect 1457 121 1463 297
rect 1417 109 1463 121
rect 1513 297 1559 309
rect 1513 121 1519 297
rect 1553 121 1559 297
rect 1513 109 1559 121
rect 1609 297 1655 309
rect 1609 121 1615 297
rect 1649 121 1655 297
rect 1609 109 1655 121
rect 1705 297 1751 309
rect 1705 121 1711 297
rect 1745 121 1751 297
rect 1705 109 1751 121
rect 1801 297 1847 309
rect 1801 121 1807 297
rect 1841 121 1847 297
rect 1801 109 1847 121
rect 1897 297 1943 309
rect 1897 121 1903 297
rect 1937 121 1943 297
rect 1897 109 1943 121
rect -1805 71 -1747 77
rect -1805 37 -1793 71
rect -1759 37 -1747 71
rect -1805 31 -1747 37
rect -1613 71 -1555 77
rect -1613 37 -1601 71
rect -1567 37 -1555 71
rect -1613 31 -1555 37
rect -1421 71 -1363 77
rect -1421 37 -1409 71
rect -1375 37 -1363 71
rect -1421 31 -1363 37
rect -1229 71 -1171 77
rect -1229 37 -1217 71
rect -1183 37 -1171 71
rect -1229 31 -1171 37
rect -1037 71 -979 77
rect -1037 37 -1025 71
rect -991 37 -979 71
rect -1037 31 -979 37
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect 1075 71 1133 77
rect 1075 37 1087 71
rect 1121 37 1133 71
rect 1075 31 1133 37
rect 1267 71 1325 77
rect 1267 37 1279 71
rect 1313 37 1325 71
rect 1267 31 1325 37
rect 1459 71 1517 77
rect 1459 37 1471 71
rect 1505 37 1517 71
rect 1459 31 1517 37
rect 1651 71 1709 77
rect 1651 37 1663 71
rect 1697 37 1709 71
rect 1651 31 1709 37
rect 1843 71 1901 77
rect 1843 37 1855 71
rect 1889 37 1901 71
rect 1843 31 1901 37
rect -1805 -37 -1747 -31
rect -1805 -71 -1793 -37
rect -1759 -71 -1747 -37
rect -1805 -77 -1747 -71
rect -1613 -37 -1555 -31
rect -1613 -71 -1601 -37
rect -1567 -71 -1555 -37
rect -1613 -77 -1555 -71
rect -1421 -37 -1363 -31
rect -1421 -71 -1409 -37
rect -1375 -71 -1363 -37
rect -1421 -77 -1363 -71
rect -1229 -37 -1171 -31
rect -1229 -71 -1217 -37
rect -1183 -71 -1171 -37
rect -1229 -77 -1171 -71
rect -1037 -37 -979 -31
rect -1037 -71 -1025 -37
rect -991 -71 -979 -37
rect -1037 -77 -979 -71
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect 1075 -37 1133 -31
rect 1075 -71 1087 -37
rect 1121 -71 1133 -37
rect 1075 -77 1133 -71
rect 1267 -37 1325 -31
rect 1267 -71 1279 -37
rect 1313 -71 1325 -37
rect 1267 -77 1325 -71
rect 1459 -37 1517 -31
rect 1459 -71 1471 -37
rect 1505 -71 1517 -37
rect 1459 -77 1517 -71
rect 1651 -37 1709 -31
rect 1651 -71 1663 -37
rect 1697 -71 1709 -37
rect 1651 -77 1709 -71
rect 1843 -37 1901 -31
rect 1843 -71 1855 -37
rect 1889 -71 1901 -37
rect 1843 -77 1901 -71
rect -1943 -121 -1897 -109
rect -1943 -297 -1937 -121
rect -1903 -297 -1897 -121
rect -1943 -309 -1897 -297
rect -1847 -121 -1801 -109
rect -1847 -297 -1841 -121
rect -1807 -297 -1801 -121
rect -1847 -309 -1801 -297
rect -1751 -121 -1705 -109
rect -1751 -297 -1745 -121
rect -1711 -297 -1705 -121
rect -1751 -309 -1705 -297
rect -1655 -121 -1609 -109
rect -1655 -297 -1649 -121
rect -1615 -297 -1609 -121
rect -1655 -309 -1609 -297
rect -1559 -121 -1513 -109
rect -1559 -297 -1553 -121
rect -1519 -297 -1513 -121
rect -1559 -309 -1513 -297
rect -1463 -121 -1417 -109
rect -1463 -297 -1457 -121
rect -1423 -297 -1417 -121
rect -1463 -309 -1417 -297
rect -1367 -121 -1321 -109
rect -1367 -297 -1361 -121
rect -1327 -297 -1321 -121
rect -1367 -309 -1321 -297
rect -1271 -121 -1225 -109
rect -1271 -297 -1265 -121
rect -1231 -297 -1225 -121
rect -1271 -309 -1225 -297
rect -1175 -121 -1129 -109
rect -1175 -297 -1169 -121
rect -1135 -297 -1129 -121
rect -1175 -309 -1129 -297
rect -1079 -121 -1033 -109
rect -1079 -297 -1073 -121
rect -1039 -297 -1033 -121
rect -1079 -309 -1033 -297
rect -983 -121 -937 -109
rect -983 -297 -977 -121
rect -943 -297 -937 -121
rect -983 -309 -937 -297
rect -887 -121 -841 -109
rect -887 -297 -881 -121
rect -847 -297 -841 -121
rect -887 -309 -841 -297
rect -791 -121 -745 -109
rect -791 -297 -785 -121
rect -751 -297 -745 -121
rect -791 -309 -745 -297
rect -695 -121 -649 -109
rect -695 -297 -689 -121
rect -655 -297 -649 -121
rect -695 -309 -649 -297
rect -599 -121 -553 -109
rect -599 -297 -593 -121
rect -559 -297 -553 -121
rect -599 -309 -553 -297
rect -503 -121 -457 -109
rect -503 -297 -497 -121
rect -463 -297 -457 -121
rect -503 -309 -457 -297
rect -407 -121 -361 -109
rect -407 -297 -401 -121
rect -367 -297 -361 -121
rect -407 -309 -361 -297
rect -311 -121 -265 -109
rect -311 -297 -305 -121
rect -271 -297 -265 -121
rect -311 -309 -265 -297
rect -215 -121 -169 -109
rect -215 -297 -209 -121
rect -175 -297 -169 -121
rect -215 -309 -169 -297
rect -119 -121 -73 -109
rect -119 -297 -113 -121
rect -79 -297 -73 -121
rect -119 -309 -73 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 73 -121 119 -109
rect 73 -297 79 -121
rect 113 -297 119 -121
rect 73 -309 119 -297
rect 169 -121 215 -109
rect 169 -297 175 -121
rect 209 -297 215 -121
rect 169 -309 215 -297
rect 265 -121 311 -109
rect 265 -297 271 -121
rect 305 -297 311 -121
rect 265 -309 311 -297
rect 361 -121 407 -109
rect 361 -297 367 -121
rect 401 -297 407 -121
rect 361 -309 407 -297
rect 457 -121 503 -109
rect 457 -297 463 -121
rect 497 -297 503 -121
rect 457 -309 503 -297
rect 553 -121 599 -109
rect 553 -297 559 -121
rect 593 -297 599 -121
rect 553 -309 599 -297
rect 649 -121 695 -109
rect 649 -297 655 -121
rect 689 -297 695 -121
rect 649 -309 695 -297
rect 745 -121 791 -109
rect 745 -297 751 -121
rect 785 -297 791 -121
rect 745 -309 791 -297
rect 841 -121 887 -109
rect 841 -297 847 -121
rect 881 -297 887 -121
rect 841 -309 887 -297
rect 937 -121 983 -109
rect 937 -297 943 -121
rect 977 -297 983 -121
rect 937 -309 983 -297
rect 1033 -121 1079 -109
rect 1033 -297 1039 -121
rect 1073 -297 1079 -121
rect 1033 -309 1079 -297
rect 1129 -121 1175 -109
rect 1129 -297 1135 -121
rect 1169 -297 1175 -121
rect 1129 -309 1175 -297
rect 1225 -121 1271 -109
rect 1225 -297 1231 -121
rect 1265 -297 1271 -121
rect 1225 -309 1271 -297
rect 1321 -121 1367 -109
rect 1321 -297 1327 -121
rect 1361 -297 1367 -121
rect 1321 -309 1367 -297
rect 1417 -121 1463 -109
rect 1417 -297 1423 -121
rect 1457 -297 1463 -121
rect 1417 -309 1463 -297
rect 1513 -121 1559 -109
rect 1513 -297 1519 -121
rect 1553 -297 1559 -121
rect 1513 -309 1559 -297
rect 1609 -121 1655 -109
rect 1609 -297 1615 -121
rect 1649 -297 1655 -121
rect 1609 -309 1655 -297
rect 1705 -121 1751 -109
rect 1705 -297 1711 -121
rect 1745 -297 1751 -121
rect 1705 -309 1751 -297
rect 1801 -121 1847 -109
rect 1801 -297 1807 -121
rect 1841 -297 1847 -121
rect 1801 -309 1847 -297
rect 1897 -121 1943 -109
rect 1897 -297 1903 -121
rect 1937 -297 1943 -121
rect 1897 -309 1943 -297
rect -1901 -347 -1843 -341
rect -1901 -381 -1889 -347
rect -1855 -381 -1843 -347
rect -1901 -387 -1843 -381
rect -1709 -347 -1651 -341
rect -1709 -381 -1697 -347
rect -1663 -381 -1651 -347
rect -1709 -387 -1651 -381
rect -1517 -347 -1459 -341
rect -1517 -381 -1505 -347
rect -1471 -381 -1459 -347
rect -1517 -387 -1459 -381
rect -1325 -347 -1267 -341
rect -1325 -381 -1313 -347
rect -1279 -381 -1267 -347
rect -1325 -387 -1267 -381
rect -1133 -347 -1075 -341
rect -1133 -381 -1121 -347
rect -1087 -381 -1075 -347
rect -1133 -387 -1075 -381
rect -941 -347 -883 -341
rect -941 -381 -929 -347
rect -895 -381 -883 -347
rect -941 -387 -883 -381
rect -749 -347 -691 -341
rect -749 -381 -737 -347
rect -703 -381 -691 -347
rect -749 -387 -691 -381
rect -557 -347 -499 -341
rect -557 -381 -545 -347
rect -511 -381 -499 -347
rect -557 -387 -499 -381
rect -365 -347 -307 -341
rect -365 -381 -353 -347
rect -319 -381 -307 -347
rect -365 -387 -307 -381
rect -173 -347 -115 -341
rect -173 -381 -161 -347
rect -127 -381 -115 -347
rect -173 -387 -115 -381
rect 19 -347 77 -341
rect 19 -381 31 -347
rect 65 -381 77 -347
rect 19 -387 77 -381
rect 211 -347 269 -341
rect 211 -381 223 -347
rect 257 -381 269 -347
rect 211 -387 269 -381
rect 403 -347 461 -341
rect 403 -381 415 -347
rect 449 -381 461 -347
rect 403 -387 461 -381
rect 595 -347 653 -341
rect 595 -381 607 -347
rect 641 -381 653 -347
rect 595 -387 653 -381
rect 787 -347 845 -341
rect 787 -381 799 -347
rect 833 -381 845 -347
rect 787 -387 845 -381
rect 979 -347 1037 -341
rect 979 -381 991 -347
rect 1025 -381 1037 -347
rect 979 -387 1037 -381
rect 1171 -347 1229 -341
rect 1171 -381 1183 -347
rect 1217 -381 1229 -347
rect 1171 -387 1229 -381
rect 1363 -347 1421 -341
rect 1363 -381 1375 -347
rect 1409 -381 1421 -347
rect 1363 -387 1421 -381
rect 1555 -347 1613 -341
rect 1555 -381 1567 -347
rect 1601 -381 1613 -347
rect 1555 -387 1613 -381
rect 1747 -347 1805 -341
rect 1747 -381 1759 -347
rect 1793 -381 1805 -347
rect 1747 -387 1805 -381
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -2034 -466 2034 466
string parameters w 1 l 0.150 m 2 nf 40 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
