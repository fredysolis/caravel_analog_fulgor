magic
tech sky130A
magscale 1 2
timestamp 1623980668
<< pwell >>
rect -16462 -24206 34360 5780
<< psubdiff >>
rect -16450 4360 -14850 4384
rect 32749 4360 34349 4384
rect 151 -145 175 -79
rect 4035 -145 4059 -79
rect -16450 -21664 -14850 -21640
rect -16450 -22594 -14851 -21664
rect 32749 -22593 34349 -21640
rect 32749 -22594 34348 -22593
rect -16450 -24194 -11039 -22594
rect 28961 -24194 34348 -22594
<< psubdiffcont >>
rect -16450 -21640 -14850 4360
rect 175 -145 4035 -79
rect 32749 -21640 34349 4360
rect -11039 -24194 28961 -22594
<< locali >>
rect -16450 4360 -14850 4376
rect 32749 4360 34349 4376
rect -14851 -21656 -14850 -21640
rect 34348 -21656 34349 -21640
<< viali >>
rect -16450 -21640 -14850 4360
rect 36 36 4230 70
rect 36 -79 4224 -49
rect 36 -145 175 -79
rect 175 -145 4035 -79
rect 4035 -145 4224 -79
rect 36 -168 4224 -145
rect -7067 -9695 -6984 -8740
rect -16450 -22594 -14851 -21640
rect 32749 -21640 34349 4360
rect 32749 -22594 34348 -21640
rect -16450 -24194 -11039 -22594
rect -11039 -24194 28961 -22594
rect 28961 -24194 34348 -22594
<< metal1 >>
rect -370 5080 -360 5680
rect 640 5614 650 5680
rect 2456 5614 2466 5680
rect 640 5182 1312 5614
rect 1560 5182 2466 5614
rect 640 5080 650 5182
rect 2456 5080 2466 5182
rect 3866 5614 3876 5680
rect 3866 5182 4100 5614
rect 3866 5080 3876 5182
rect -16456 4360 -14844 4372
rect -16456 -21634 -16450 4360
rect -16462 -24194 -16450 -21634
rect -14850 -21634 -14844 4360
rect 32743 4360 34355 4372
rect 166 166 3245 598
rect -10 70 4297 90
rect -10 36 36 70
rect 4230 36 4297 70
rect -10 -49 4297 36
rect -10 -168 36 -49
rect 4224 -168 4297 -49
rect -10 -185 4297 -168
rect 1312 -1221 2954 -185
rect 1312 -1273 2955 -1221
rect 1313 -2326 2955 -1273
rect -7073 -8740 -6978 -8728
rect -7325 -9502 -7315 -8929
rect -7258 -9502 -7248 -8929
rect -7191 -9505 -7181 -8922
rect -7129 -9505 -7119 -8922
rect -7073 -9695 -7067 -8740
rect -6984 -8828 -6978 -8740
rect -6903 -9581 -6893 -8828
rect -6984 -9695 -6978 -9581
rect -7073 -9707 -6978 -9695
rect -14850 -21640 -14839 -21634
rect -14851 -22588 -14839 -21640
rect 1313 -22588 2954 -2326
rect 32743 -22588 32749 4360
rect 34349 -21640 34355 4360
rect -14851 -22594 32749 -22588
rect 34348 -21652 34355 -21640
rect 34348 -22588 34354 -21652
rect 34348 -24194 34360 -22588
rect -16462 -24200 34360 -24194
rect 32743 -24206 34354 -24200
<< via1 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -7315 -9502 -7258 -8929
rect -7181 -9505 -7129 -8922
rect -7009 -9581 -6984 -8828
rect -6984 -9581 -6903 -8828
rect -10029 -23953 -4329 -22753
rect 9433 -24034 31413 -22834
<< metal2 >>
rect -360 5680 640 5690
rect -360 5070 640 5080
rect 2466 5680 3866 5690
rect 2466 5070 3866 5080
rect -6973 -8818 -6867 -8814
rect -7009 -8824 -6867 -8818
rect -7009 -8828 -6973 -8824
rect -7181 -8913 -7129 -8912
rect -7315 -8920 -7258 -8919
rect -7334 -8929 -7258 -8920
rect -7334 -8930 -7315 -8929
rect -7267 -9503 -7258 -9502
rect -7334 -9512 -7258 -9503
rect -7181 -8922 -7114 -8913
rect -7129 -8923 -7114 -8922
rect -7334 -9513 -7267 -9512
rect -7181 -9515 -7114 -9505
rect -6903 -9581 -6867 -9577
rect -7009 -9587 -6867 -9581
rect -7009 -9591 -6903 -9587
rect -10029 -22753 -4329 -22743
rect -10029 -23963 -4329 -23953
rect 9433 -22834 31413 -22824
rect 9433 -24044 31413 -24034
<< via2 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -6973 -8828 -6867 -8824
rect -7334 -9502 -7315 -8930
rect -7315 -9502 -7267 -8930
rect -7334 -9503 -7267 -9502
rect -7181 -9505 -7129 -8923
rect -7129 -9505 -7114 -8923
rect -6973 -9577 -6903 -8828
rect -6903 -9577 -6867 -8828
rect -10029 -23953 -4329 -22753
rect 9433 -24034 31413 -22834
<< metal3 >>
rect -370 5680 650 5685
rect -370 5080 -360 5680
rect 640 5080 650 5680
rect -370 5075 650 5080
rect 2456 5680 3876 5685
rect 2456 5080 2466 5680
rect 3866 5080 3876 5680
rect 2456 5075 3876 5080
rect -13523 -8002 -586 4898
rect -10029 -10424 -8629 -8002
rect -6983 -8824 -6857 -8819
rect -7191 -8923 -7104 -8918
rect -7344 -8928 -7257 -8925
rect -7379 -9504 -7369 -8928
rect -7264 -9504 -7254 -8928
rect -7344 -9508 -7257 -9504
rect -7191 -9505 -7181 -8923
rect -7082 -9505 -7072 -8923
rect -7191 -9510 -7104 -9505
rect -6983 -9577 -6973 -8824
rect -6867 -8830 -6857 -8824
rect -5695 -8830 -4295 -8002
rect -6867 -9577 -4295 -8830
rect -6983 -9582 -6857 -9577
rect -5695 -10424 -4295 -9577
rect -11511 -19024 -2893 -10424
rect -10029 -22748 -8629 -19024
rect -5695 -22748 -4295 -19024
rect 4852 -21602 31427 4898
rect -10039 -22753 -4295 -22748
rect -10039 -23953 -10029 -22753
rect -4329 -23136 -4295 -22753
rect 9433 -22829 10833 -21602
rect 14842 -22829 16242 -21602
rect 20055 -22829 21455 -21602
rect 25394 -22829 26794 -21602
rect 30027 -22829 31427 -21602
rect 9423 -22834 31427 -22829
rect -4329 -23953 -4319 -23136
rect -10039 -23958 -4319 -23953
rect 9423 -24034 9433 -22834
rect 31413 -23602 31427 -22834
rect 31413 -24034 31423 -23602
rect 9423 -24039 31423 -24034
rect 25394 -24061 26794 -24039
<< via3 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -7369 -8930 -7264 -8928
rect -7369 -9503 -7334 -8930
rect -7334 -9503 -7267 -8930
rect -7267 -9503 -7264 -8930
rect -7369 -9504 -7264 -9503
rect -7181 -9505 -7114 -8923
rect -7114 -9505 -7082 -8923
<< metal4 >>
rect -12154 5680 740 5780
rect -12154 5080 -360 5680
rect 640 5080 740 5680
rect -12154 4980 740 5080
rect 2066 5680 29520 5780
rect 2066 5080 2466 5680
rect 3866 5080 29520 5680
rect 2066 4980 29520 5080
rect -12154 -6696 -10754 4980
rect -7779 -6696 -6379 4980
rect -3405 -6534 -2005 4980
rect -11475 -8112 -11371 -7898
rect -7156 -8112 -7052 -7866
rect -2837 -8112 -2733 -7848
rect -11475 -8216 -2733 -8112
rect -7369 -8927 -7263 -8216
rect -7182 -8923 -7081 -8922
rect -7182 -8924 -7181 -8923
rect -7370 -8928 -7263 -8927
rect -7370 -9504 -7369 -8928
rect -7264 -9504 -7263 -8928
rect -7370 -9505 -7263 -9504
rect -7183 -9505 -7181 -8924
rect -7082 -8924 -7081 -8923
rect -7082 -9505 -7077 -8924
rect -7183 -10154 -7077 -9505
rect -9463 -10258 -5040 -10154
rect -9463 -10536 -9359 -10258
rect -5144 -10528 -5040 -10258
rect -9463 -19216 -9359 -18920
rect -5144 -19216 -5040 -18920
rect 6722 -19031 8122 4980
rect 12166 -19023 13566 4980
rect 17484 -19174 18884 4980
rect -9463 -19320 -5040 -19216
rect 22862 -19265 24262 4980
rect 28119 -19235 29519 4980
rect -5144 -19321 -5040 -19320
use sky130_fd_pr__nfet_01v8_U2JGXT  sky130_fd_pr__nfet_01v8_U2JGXT_0
timestamp 1623980668
transform 1 0 -7220 0 1 -9214
box -226 -510 226 510
use sky130_fd_pr__cap_mim_m3_1_BC3K5K  sky130_fd_pr__cap_mim_m3_1_BC3K5K_0
timestamp 1623980668
transform 1 0 -7202 0 1 -14724
box -4309 -4300 4309 4300
use sky130_fd_pr__res_high_po_5p73_GW5RGE  sky130_fd_pr__res_high_po_5p73_GW5RGE_0
timestamp 1623892191
transform 1 0 2133 0 1 2890
box -2133 -2890 2133 2890
use sky130_fd_pr__cap_mim_m3_1_MA89VW  sky130_fd_pr__cap_mim_m3_1_MA89VW_0
timestamp 1623892191
transform 1 0 18140 0 1 -8352
box -13288 -13250 13287 13250
use sky130_fd_pr__cap_mim_m3_1_W3JTNJ  sky130_fd_pr__cap_mim_m3_1_W3JTNJ_0
timestamp 1623892191
transform 1 0 -7054 0 1 -1552
box -6469 -6450 6468 6450
<< labels >>
rlabel metal4 3866 4980 29520 5780 1 vc_pex
rlabel metal4 -12154 4980 -360 5780 1 in
rlabel metal1 1313 -22594 2954 -168 1 vss
<< end >>
