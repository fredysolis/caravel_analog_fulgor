magic
tech sky130A
magscale 1 2
timestamp 1623943772
<< error_p >>
rect -173 385 -115 391
rect 19 385 77 391
rect -173 351 -161 385
rect 19 351 31 385
rect -173 345 -115 351
rect 19 345 77 351
rect -77 71 -19 77
rect 115 71 173 77
rect -77 37 -65 71
rect 115 37 127 71
rect -77 31 -19 37
rect 115 31 173 37
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect -173 -351 -115 -345
rect 19 -351 77 -345
rect -173 -385 -161 -351
rect 19 -385 31 -351
rect -173 -391 -115 -385
rect 19 -391 77 -385
<< pwell >>
rect -359 -523 359 523
<< nmos >>
rect -159 109 -129 313
rect -63 109 -33 313
rect 33 109 63 313
rect 129 109 159 313
rect -159 -313 -129 -109
rect -63 -313 -33 -109
rect 33 -313 63 -109
rect 129 -313 159 -109
<< ndiff >>
rect -221 301 -159 313
rect -221 121 -209 301
rect -175 121 -159 301
rect -221 109 -159 121
rect -129 301 -63 313
rect -129 121 -113 301
rect -79 121 -63 301
rect -129 109 -63 121
rect -33 301 33 313
rect -33 121 -17 301
rect 17 121 33 301
rect -33 109 33 121
rect 63 301 129 313
rect 63 121 79 301
rect 113 121 129 301
rect 63 109 129 121
rect 159 301 221 313
rect 159 121 175 301
rect 209 121 221 301
rect 159 109 221 121
rect -221 -121 -159 -109
rect -221 -301 -209 -121
rect -175 -301 -159 -121
rect -221 -313 -159 -301
rect -129 -121 -63 -109
rect -129 -301 -113 -121
rect -79 -301 -63 -121
rect -129 -313 -63 -301
rect -33 -121 33 -109
rect -33 -301 -17 -121
rect 17 -301 33 -121
rect -33 -313 33 -301
rect 63 -121 129 -109
rect 63 -301 79 -121
rect 113 -301 129 -121
rect 63 -313 129 -301
rect 159 -121 221 -109
rect 159 -301 175 -121
rect 209 -301 221 -121
rect 159 -313 221 -301
<< ndiffc >>
rect -209 121 -175 301
rect -113 121 -79 301
rect -17 121 17 301
rect 79 121 113 301
rect 175 121 209 301
rect -209 -301 -175 -121
rect -113 -301 -79 -121
rect -17 -301 17 -121
rect 79 -301 113 -121
rect 175 -301 209 -121
<< psubdiff >>
rect -323 453 323 487
rect -323 391 -289 453
rect 289 391 323 453
rect -323 -453 -289 -391
rect 289 -453 323 -391
rect -323 -487 -227 -453
rect 227 -487 323 -453
<< psubdiffcont >>
rect -323 -391 -289 391
rect 289 -391 323 391
rect -227 -487 227 -453
<< poly >>
rect -177 385 -111 401
rect -177 351 -161 385
rect -127 351 -111 385
rect -177 335 -111 351
rect 15 385 81 401
rect 15 351 31 385
rect 65 351 81 385
rect -159 313 -129 335
rect -63 313 -33 339
rect 15 335 81 351
rect 33 313 63 335
rect 129 313 159 339
rect -159 83 -129 109
rect -63 87 -33 109
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 129 -109 159 -87
rect -159 -335 -129 -313
rect -177 -351 -111 -335
rect -63 -339 -33 -313
rect 33 -335 63 -313
rect -177 -385 -161 -351
rect -127 -385 -111 -351
rect -177 -401 -111 -385
rect 15 -351 81 -335
rect 129 -339 159 -313
rect 15 -385 31 -351
rect 65 -385 81 -351
rect 15 -401 81 -385
<< polycont >>
rect -161 351 -127 385
rect 31 351 65 385
rect -65 37 -31 71
rect 127 37 161 71
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect -161 -385 -127 -351
rect 31 -385 65 -351
<< locali >>
rect -323 453 323 487
rect -323 391 -289 453
rect 289 391 323 453
rect -177 351 -161 385
rect -127 351 -111 385
rect 15 351 31 385
rect 65 351 81 385
rect -209 301 -175 317
rect -209 105 -175 121
rect -113 301 -79 317
rect -113 105 -79 121
rect -17 301 17 317
rect -17 105 17 121
rect 79 301 113 317
rect 79 105 113 121
rect 175 301 209 317
rect 175 105 209 121
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -209 -121 -175 -105
rect -209 -317 -175 -301
rect -113 -121 -79 -105
rect -113 -317 -79 -301
rect -17 -121 17 -105
rect -17 -317 17 -301
rect 79 -121 113 -105
rect 79 -317 113 -301
rect 175 -121 209 -105
rect 175 -317 209 -301
rect -177 -385 -161 -351
rect -127 -385 -111 -351
rect 15 -385 31 -351
rect 65 -385 81 -351
rect -323 -453 -289 -391
rect 289 -453 323 -391
rect -323 -487 -227 -453
rect 227 -487 323 -453
<< viali >>
rect -161 351 -127 385
rect 31 351 65 385
rect -209 121 -175 301
rect -113 121 -79 301
rect -17 121 17 301
rect 79 121 113 301
rect 175 121 209 301
rect -65 37 -31 71
rect 127 37 161 71
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect -209 -301 -175 -121
rect -113 -301 -79 -121
rect -17 -301 17 -121
rect 79 -301 113 -121
rect 175 -301 209 -121
rect -161 -385 -127 -351
rect 31 -385 65 -351
<< metal1 >>
rect -173 385 -115 391
rect -173 351 -161 385
rect -127 351 -115 385
rect -173 345 -115 351
rect 19 385 77 391
rect 19 351 31 385
rect 65 351 77 385
rect 19 345 77 351
rect -215 301 -169 313
rect -215 121 -209 301
rect -175 121 -169 301
rect -215 109 -169 121
rect -119 301 -73 313
rect -119 121 -113 301
rect -79 121 -73 301
rect -119 109 -73 121
rect -23 301 23 313
rect -23 121 -17 301
rect 17 121 23 301
rect -23 109 23 121
rect 73 301 119 313
rect 73 121 79 301
rect 113 121 119 301
rect 73 109 119 121
rect 169 301 215 313
rect 169 121 175 301
rect 209 121 215 301
rect 169 109 215 121
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect -215 -121 -169 -109
rect -215 -301 -209 -121
rect -175 -301 -169 -121
rect -215 -313 -169 -301
rect -119 -121 -73 -109
rect -119 -301 -113 -121
rect -79 -301 -73 -121
rect -119 -313 -73 -301
rect -23 -121 23 -109
rect -23 -301 -17 -121
rect 17 -301 23 -121
rect -23 -313 23 -301
rect 73 -121 119 -109
rect 73 -301 79 -121
rect 113 -301 119 -121
rect 73 -313 119 -301
rect 169 -121 215 -109
rect 169 -301 175 -121
rect 209 -301 215 -121
rect 169 -313 215 -301
rect -173 -351 -115 -345
rect -173 -385 -161 -351
rect -127 -385 -115 -351
rect -173 -391 -115 -385
rect 19 -351 77 -345
rect 19 -385 31 -351
rect 65 -385 77 -351
rect 19 -391 77 -385
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -306 -470 306 470
string parameters w 1.02 l 0.150 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
