magic
tech sky130A
magscale 1 2
timestamp 1624046389
<< nwell >>
rect -53 531 1817 643
rect -31 -19 1817 531
rect -31 -53 574 -19
rect 1037 -53 1817 -19
<< pwell >>
rect -18 -610 1781 -576
<< psubdiff >>
rect -17 -610 79 -576
rect 1685 -610 1781 -576
<< nsubdiff >>
rect -17 571 79 605
rect 1685 571 1781 605
<< psubdiffcont >>
rect 79 -610 1685 -576
<< nsubdiffcont >>
rect 79 571 1685 605
<< poly >>
rect 147 83 465 140
rect 147 81 300 83
rect 147 10 930 81
rect 147 -123 190 10
rect 258 -123 930 10
rect 147 -175 930 -123
rect 147 -181 300 -175
rect 147 -238 465 -181
<< polycont >>
rect 190 -123 258 10
<< locali >>
rect 174 10 274 26
rect 174 -123 190 10
rect 258 -123 274 10
rect 174 -139 274 -123
<< viali >>
rect -17 571 79 605
rect 79 571 1685 605
rect 1685 571 1782 605
rect -17 483 1782 517
rect 190 -123 258 10
rect -18 -521 1781 -487
rect -18 -610 79 -576
rect 79 -610 1685 -576
rect 1685 -610 1781 -576
<< metal1 >>
rect 665 611 1817 612
rect -53 605 1817 611
rect -53 571 -17 605
rect 1782 571 1817 605
rect -53 517 1817 571
rect -53 483 -17 517
rect 1782 483 1817 517
rect -53 477 1817 483
rect 88 129 137 334
rect 177 166 243 477
rect 281 129 330 333
rect 369 166 435 477
rect 475 129 521 185
rect 561 166 627 477
rect 667 129 713 190
rect 753 166 819 477
rect 859 129 905 188
rect 945 166 1011 477
rect 1051 129 1097 187
rect 1137 166 1203 477
rect 1243 129 1289 187
rect 1329 166 1395 477
rect 1435 129 1481 188
rect 1521 166 1587 477
rect 1627 129 1673 184
rect 88 59 1675 129
rect 184 10 264 22
rect 184 -13 190 10
rect -53 -93 190 -13
rect 184 -123 190 -93
rect 258 -123 264 10
rect 184 -135 264 -123
rect 1034 -19 1675 59
rect 1034 -97 1817 -19
rect 1034 -165 1675 -97
rect 90 -232 1675 -165
rect 90 -347 139 -232
rect 177 -481 243 -262
rect 282 -348 331 -232
rect 369 -481 435 -261
rect 475 -283 521 -232
rect 561 -481 627 -261
rect 667 -276 713 -232
rect 753 -481 819 -261
rect 859 -272 905 -232
rect 945 -481 1011 -263
rect 1051 -273 1097 -232
rect 1137 -481 1203 -263
rect 1243 -273 1289 -232
rect 1329 -481 1395 -263
rect 1435 -271 1481 -232
rect 1521 -481 1587 -263
rect 1627 -270 1673 -232
rect -53 -487 1817 -481
rect -53 -521 -18 -487
rect 1781 -521 1817 -487
rect -53 -576 1817 -521
rect -53 -610 -18 -576
rect 1781 -610 1817 -576
rect -53 -616 1817 -610
use sky130_fd_pr__pfet_01v8_BDRUME  sky130_fd_pr__pfet_01v8_BDRUME_0
timestamp 1624046389
transform 1 0 882 0 1 250
box -935 -303 935 303
use sky130_fd_pr__nfet_01v8_QQE8KM  sky130_fd_pr__nfet_01v8_QQE8KM_0
timestamp 1624046389
transform 1 0 882 0 1 -305
box -935 -252 935 252
<< labels >>
rlabel metal1 -53 -576 665 -521 1 vss
rlabel metal1 -53 -93 190 -13 1 in
rlabel metal1 -53 517 665 571 1 vdd
rlabel metal1 1650 -97 1817 -19 1 out
<< end >>
