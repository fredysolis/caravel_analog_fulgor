magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect -422 2867 0 2956
<< pwell >>
rect 1294 809 1725 1389
rect 2588 809 3019 1389
rect -422 165 -411 166
rect -422 0 0 165
<< psubdiff >>
rect -314 36 -290 70
rect -132 36 -108 70
<< nsubdiff >>
rect -314 2886 -290 2920
rect -132 2886 -108 2920
<< psubdiffcont >>
rect -290 36 -132 70
<< nsubdiffcont >>
rect -290 2886 -132 2920
<< viali >>
rect -386 2886 -290 2920
rect -290 2886 -132 2920
rect -132 2886 -36 2920
rect -386 2797 -36 2831
rect -386 125 -36 159
rect -386 36 -290 70
rect -290 36 -132 70
rect -132 36 -36 70
<< metal1 >>
rect -422 2920 0 2926
rect -422 2886 -386 2920
rect -36 2886 0 2920
rect -422 2831 0 2886
rect -422 2797 -386 2831
rect -36 2797 0 2831
rect -422 2791 0 2797
rect -324 2348 -278 2791
rect -243 2695 -233 2747
rect -129 2695 -119 2747
rect -243 2686 -144 2695
rect -190 2646 -144 2686
rect -190 2199 -144 2353
rect -236 739 -98 2199
rect 1294 779 1725 957
rect 2588 779 3019 957
rect -324 165 -278 599
rect -190 597 -144 739
rect -243 261 -119 270
rect -243 209 -233 261
rect -129 209 -119 261
rect -422 159 0 165
rect -422 125 -386 159
rect -36 125 0 159
rect -422 70 0 125
rect -422 36 -386 70
rect -36 36 0 70
rect -422 30 0 36
<< via1 >>
rect -233 2695 -129 2747
rect -233 209 -129 261
<< metal2 >>
rect -233 2747 3061 2757
rect -129 2695 3061 2747
rect -233 2685 3061 2695
rect 440 1417 608 1427
rect 3316 1417 3440 1427
rect 1255 1363 1757 1415
rect 2557 1363 3030 1415
rect 440 1351 608 1361
rect 3651 1363 3882 1415
rect 3316 1351 3440 1361
rect -233 261 2860 271
rect -129 209 2860 261
rect -233 199 2860 209
rect 1015 159 1071 169
rect 2309 159 2365 169
rect 3603 159 3659 169
rect 1005 103 1015 159
rect 1071 103 2309 159
rect 2365 103 3603 159
rect 3659 103 3669 159
rect 1015 94 1071 103
rect 2309 94 2365 103
rect 3603 94 3659 103
<< via2 >>
rect 440 1361 608 1417
rect 3316 1361 3440 1417
rect 1015 103 1071 159
rect 2309 103 2365 159
rect 3603 103 3659 159
<< metal3 >>
rect 430 1421 618 1422
rect 430 1417 441 1421
rect 607 1417 618 1421
rect 430 1361 440 1417
rect 608 1361 618 1417
rect 430 1357 441 1361
rect 607 1357 618 1361
rect 430 1356 618 1357
rect 3306 1421 3450 1425
rect 3306 1417 3317 1421
rect 3306 1361 3316 1417
rect 3306 1357 3317 1361
rect 3440 1357 3450 1421
rect 3306 1353 3450 1357
rect 1013 164 1073 970
rect 2307 164 2367 1007
rect 3601 164 3661 1007
rect 1005 159 1081 164
rect 1005 103 1015 159
rect 1071 103 1081 159
rect 1005 98 1081 103
rect 2299 159 2375 164
rect 2299 103 2309 159
rect 2365 103 2375 159
rect 2299 98 2375 103
rect 3593 159 3669 164
rect 3593 103 3603 159
rect 3659 103 3669 159
rect 3593 98 3669 103
rect 1013 94 1073 98
rect 2307 90 2367 98
<< via3 >>
rect 441 1417 607 1421
rect 441 1361 607 1417
rect 441 1357 607 1361
rect 3317 1417 3440 1421
rect 3317 1361 3440 1417
rect 3317 1357 3440 1361
<< metal4 >>
rect 440 1421 608 1422
rect 3316 1421 3441 1422
rect 440 1357 441 1421
rect 607 1357 3317 1421
rect 3440 1357 3441 1421
rect 440 1356 608 1357
rect 3316 1356 3441 1357
use csvco_branch  csvco_branch_2
timestamp 1624049879
transform 1 0 2951 0 1 1002
box -363 -1002 931 1954
use csvco_branch  csvco_branch_1
timestamp 1624049879
transform 1 0 1657 0 1 1002
box -363 -1002 931 1954
use csvco_branch  csvco_branch_0
timestamp 1624049879
transform 1 0 363 0 1 1002
box -363 -1002 931 1954
use sky130_fd_pr__pfet_01v8_4757AC  sky130_fd_pr__pfet_01v8_4757AC_0
timestamp 1624049879
transform 1 0 -211 0 1 2498
box -211 -369 211 369
use sky130_fd_pr__nfet_01v8_CBAU6Y  sky130_fd_pr__nfet_01v8_CBAU6Y_0
timestamp 1624049879
transform 1 0 -211 0 1 449
box -211 -360 211 360
<< labels >>
rlabel metal2 -77 211 -25 263 1 vctrl
rlabel metal1 -422 70 0 125 1 vss
rlabel metal1 -422 2831 0 2886 1 vdd
rlabel metal2 3651 1363 3882 1415 1 out_vco
rlabel via2 2309 103 2365 159 1 D0
<< end >>
