magic
tech sky130A
magscale 1 2
timestamp 1623427697
<< pwell >>
rect -263 -64 263 252
rect -263 -66 -81 -64
rect -63 -66 -33 -64
rect -15 -66 263 -64
rect -263 -252 263 -66
<< nmos >>
rect -63 -42 -33 42
rect 33 -42 63 42
<< ndiff >>
rect -125 30 -63 42
rect -125 -30 -113 30
rect -79 -30 -63 30
rect -125 -42 -63 -30
rect -33 30 33 42
rect -33 -30 -17 30
rect 17 -30 33 30
rect -33 -42 33 -30
rect 63 30 125 42
rect 63 -30 79 30
rect 113 -30 125 30
rect 63 -42 125 -30
<< ndiffc >>
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
<< psubdiff >>
rect -227 120 -193 182
rect 193 120 227 182
rect -227 -182 -193 -120
rect 193 -182 227 -120
rect -227 -216 -131 -182
rect 131 -216 227 -182
<< psubdiffcont >>
rect -227 -120 -193 120
rect 193 -120 227 120
rect -131 -216 131 -182
<< poly >>
rect -63 42 -33 68
rect 33 42 63 68
rect -63 -68 -33 -42
rect 33 -68 63 -42
<< locali >>
rect -227 120 -193 182
rect 193 120 227 182
rect -113 30 -79 46
rect -113 -46 -79 -30
rect -17 30 17 46
rect -17 -46 17 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect -227 -182 -193 -120
rect 193 -182 227 -120
rect -227 -216 -131 -182
rect 131 -216 227 -182
<< viali >>
rect -113 -30 -79 30
rect -17 -30 17 30
rect 79 -30 113 30
<< metal1 >>
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect -23 30 23 42
rect -23 -30 -17 30
rect 17 -30 23 30
rect -23 -42 23 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -210 -199 210 199
string parameters w 0.420 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
