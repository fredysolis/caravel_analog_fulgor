* NGSPICE file created from csvco_branch_v2.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_CBSTVW a_n73_n119# a_n33_n207# w_n211_n329# a_15_n119#
X0 a_15_n119# a_n33_n207# a_n73_n119# w_n211_n329# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n73_n119# a_n33_n207# 0.02fF
C1 a_n33_n207# a_15_n119# 0.02fF
C2 a_n73_n119# a_15_n119# 0.51fF
C3 a_15_n119# w_n211_n329# 0.24fF
C4 a_n73_n119# w_n211_n329# 0.24fF
C5 a_n33_n207# w_n211_n329# 0.17fF
.ends

.subckt sky130_fd_pr__pfet_01v8_MJP3BN VSUBS a_15_n186# w_n211_n334# a_n33_145# a_n73_n186#
X0 a_15_n186# a_n33_145# a_n73_n186# w_n211_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n73_n186# a_15_n186# 0.51fF
C1 a_n73_n186# a_n33_145# 0.01fF
C2 w_n211_n334# a_15_n186# 0.21fF
C3 w_n211_n334# a_n33_145# 0.05fF
C4 w_n211_n334# a_n73_n186# 0.21fF
C5 a_15_n186# a_n33_145# 0.01fF
C6 a_15_n186# VSUBS 0.03fF
C7 a_n73_n186# VSUBS 0.03fF
C8 a_n33_145# VSUBS 0.12fF
C9 w_n211_n334# VSUBS 1.81fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EDT3AT a_15_n11# a_n33_n99# w_n211_n221# a_n73_n11#
X0 a_15_n11# a_n33_n99# a_n73_n11# w_n211_n221# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_15_n11# a_n73_n11# 0.15fF
C1 a_n33_n99# a_n73_n11# 0.02fF
C2 a_n33_n99# a_15_n11# 0.02fF
C3 a_15_n11# w_n211_n221# 0.09fF
C4 a_n73_n11# w_n211_n221# 0.09fF
C5 a_n33_n99# w_n211_n221# 0.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AQR2CW a_n33_66# a_n78_n106# w_n216_n254# a_20_n106#
X0 a_20_n106# a_n33_66# a_n78_n106# w_n216_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=200000u
C0 a_20_n106# a_n78_n106# 0.21fF
C1 a_20_n106# w_n216_n254# 0.14fF
C2 a_n78_n106# w_n216_n254# 0.14fF
C3 a_n33_66# w_n216_n254# 0.12fF
.ends

.subckt sky130_fd_pr__pfet_01v8_HRYSXS VSUBS a_n33_n211# a_n78_n114# w_n216_n334#
+ a_20_n114#
X0 a_20_n114# a_n33_n211# a_n78_n114# w_n216_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=200000u
C0 a_n78_n114# a_20_n114# 0.42fF
C1 w_n216_n334# a_20_n114# 0.20fF
C2 w_n216_n334# a_n78_n114# 0.20fF
C3 a_20_n114# VSUBS 0.03fF
C4 a_n78_n114# VSUBS 0.03fF
C5 a_n33_n211# VSUBS 0.12fF
C6 w_n216_n334# VSUBS 1.66fF
.ends

.subckt inverter_csvco in vbulkn out vbulkp vdd vss
Xsky130_fd_pr__nfet_01v8_AQR2CW_0 in vss vbulkn out sky130_fd_pr__nfet_01v8_AQR2CW
Xsky130_fd_pr__pfet_01v8_HRYSXS_0 vbulkn in vdd vbulkp out sky130_fd_pr__pfet_01v8_HRYSXS
C0 vdd vbulkp 0.04fF
C1 out in 0.11fF
C2 out vbulkp 0.08fF
C3 in vdd 0.01fF
C4 in vss 0.01fF
C5 vbulkp vbulkn 2.49fF
C6 out vbulkn 0.60fF
C7 vdd vbulkn 0.06fF
C8 in vbulkn 0.54fF
C9 vss vbulkn 0.17fF
.ends


* Top level circuit csvco_branch_v2

Xsky130_fd_pr__nfet_01v8_CBSTVW_0 inverter_csvco_0/vss vctrl vss vss sky130_fd_pr__nfet_01v8_CBSTVW
Xsky130_fd_pr__pfet_01v8_MJP3BN_0 vss vdd vdd m1_185_1641# inverter_csvco_0/vdd sky130_fd_pr__pfet_01v8_MJP3BN
Xsky130_fd_pr__nfet_01v8_EDT3AT_0 cap_vco_0/t D0 vss out sky130_fd_pr__nfet_01v8_EDT3AT
Xinverter_csvco_0 in vss out vdd inverter_csvco_0/vdd inverter_csvco_0/vss inverter_csvco
C0 inverter_csvco_0/vdd m1_185_1641# 0.13fF
C1 vdd cap_vco_0/t 0.06fF
C2 inverter_csvco_0/vss vctrl 0.23fF
C3 inverter_csvco_0/vdd cap_vco_0/t 0.10fF
C4 inverter_csvco_0/vss in 0.01fF
C5 inverter_csvco_0/vdd vdd 0.97fF
C6 inverter_csvco_0/vss out 0.03fF
C7 out cap_vco_0/t 0.70fF
C8 D0 out 0.09fF
C9 out vdd 0.03fF
C10 inverter_csvco_0/vdd in 0.01fF
C11 inverter_csvco_0/vdd out 0.02fF
C12 out in 0.06fF
C13 m1_185_1641# vdd 0.48fF
C14 inverter_csvco_0/vss D0 0.01fF
C15 vdd vss 3.61fF
C16 out vss 0.94fF
C17 inverter_csvco_0/vdd vss 0.23fF
C18 in vss 0.70fF
C19 inverter_csvco_0/vss vss 0.61fF
C20 D0 vss -0.68fF
C21 m1_185_1641# vss -0.03fF
C22 cap_vco_0/t vss 7.22fF
C23 vctrl vss 0.44fF
.end

