magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< metal3 >>
rect -8638 -8650 4299 4250
rect -7038 -8892 -6038 -8650
rect -2719 -8892 -1719 -8650
rect 1600 -8892 2600 -8650
rect -7038 -9892 2600 -8892
<< metal4 >>
rect -7038 4492 2600 5492
rect -7038 2599 -6038 4492
rect -2719 2599 -1719 4492
rect 1600 2599 2600 4492
rect -7038 1599 2600 2599
rect -7038 -1700 -6038 1599
rect -2719 -1700 -1719 1599
rect 1600 -1700 2600 1599
rect -7038 -2700 2600 -1700
rect -7038 -6000 -6038 -2700
rect -2719 -6000 -1719 -2700
rect 1600 -6000 2600 -2700
rect -7038 -7000 2600 -6000
rect -7038 -8650 -6038 -7000
rect -2719 -8650 -1719 -7000
rect 1600 -8650 2600 -7000
use sky130_fd_pr__cap_mim_m3_1_W3JTNJ  sky130_fd_pr__cap_mim_m3_1_W3JTNJ_0
timestamp 1624049879
transform 1 0 -2169 0 1 -2200
box -6469 -6450 6468 6450
<< labels >>
rlabel metal4 -7038 4492 2600 5492 1 in
rlabel metal3 -7038 -9892 2600 -8892 1 out
<< end >>
