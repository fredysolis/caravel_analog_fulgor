magic
tech sky130A
magscale 1 2
timestamp 1623947031
<< error_p >>
rect -239 181 -181 187
rect 181 181 239 187
rect -239 147 -227 181
rect 181 147 193 181
rect -239 141 -181 147
rect 181 141 239 147
rect -449 -147 -391 -141
rect -29 -147 29 -141
rect 391 -147 449 -141
rect -449 -181 -437 -147
rect -29 -181 -17 -147
rect 391 -181 403 -147
rect -449 -187 -391 -181
rect -29 -187 29 -181
rect 391 -187 449 -181
<< nwell >>
rect -635 -319 635 319
<< pmos >>
rect -435 -100 -405 100
rect -225 -100 -195 100
rect -15 -100 15 100
rect 195 -100 225 100
rect 405 -100 435 100
<< pdiff >>
rect -497 88 -435 100
rect -497 -88 -485 88
rect -451 -88 -435 88
rect -497 -100 -435 -88
rect -405 88 -343 100
rect -405 -88 -389 88
rect -355 -88 -343 88
rect -405 -100 -343 -88
rect -287 88 -225 100
rect -287 -88 -275 88
rect -241 -88 -225 88
rect -287 -100 -225 -88
rect -195 88 -133 100
rect -195 -88 -179 88
rect -145 -88 -133 88
rect -195 -100 -133 -88
rect -77 88 -15 100
rect -77 -88 -65 88
rect -31 -88 -15 88
rect -77 -100 -15 -88
rect 15 88 77 100
rect 15 -88 31 88
rect 65 -88 77 88
rect 15 -100 77 -88
rect 133 88 195 100
rect 133 -88 145 88
rect 179 -88 195 88
rect 133 -100 195 -88
rect 225 88 287 100
rect 225 -88 241 88
rect 275 -88 287 88
rect 225 -100 287 -88
rect 343 88 405 100
rect 343 -88 355 88
rect 389 -88 405 88
rect 343 -100 405 -88
rect 435 88 497 100
rect 435 -88 451 88
rect 485 -88 497 88
rect 435 -100 497 -88
<< pdiffc >>
rect -485 -88 -451 88
rect -389 -88 -355 88
rect -275 -88 -241 88
rect -179 -88 -145 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 145 -88 179 88
rect 241 -88 275 88
rect 355 -88 389 88
rect 451 -88 485 88
<< nsubdiff >>
rect -599 249 -503 283
rect 503 249 599 283
rect -599 187 -565 249
rect 565 187 599 249
rect -599 -249 -565 -187
rect 565 -249 599 -187
rect -599 -283 -503 -249
rect 503 -283 599 -249
<< nsubdiffcont >>
rect -503 249 503 283
rect -599 -187 -565 187
rect 565 -187 599 187
rect -503 -283 503 -249
<< poly >>
rect -243 181 -177 197
rect -243 147 -227 181
rect -193 147 -177 181
rect -243 131 -177 147
rect 177 181 243 197
rect 177 147 193 181
rect 227 147 243 181
rect 177 131 243 147
rect -435 100 -405 126
rect -225 100 -195 131
rect -15 100 15 126
rect 195 100 225 131
rect 405 100 435 126
rect -435 -131 -405 -100
rect -225 -126 -195 -100
rect -15 -131 15 -100
rect 195 -126 225 -100
rect 405 -131 435 -100
rect -453 -147 -387 -131
rect -453 -181 -437 -147
rect -403 -181 -387 -147
rect -453 -197 -387 -181
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
rect 387 -147 453 -131
rect 387 -181 403 -147
rect 437 -181 453 -147
rect 387 -197 453 -181
<< polycont >>
rect -227 147 -193 181
rect 193 147 227 181
rect -437 -181 -403 -147
rect -17 -181 17 -147
rect 403 -181 437 -147
<< locali >>
rect -599 249 -503 283
rect 503 249 599 283
rect -599 187 -565 249
rect 565 187 599 249
rect -243 147 -227 181
rect -193 147 -177 181
rect 177 147 193 181
rect 227 147 243 181
rect -485 88 -451 104
rect -485 -104 -451 -88
rect -389 88 -355 104
rect -389 -104 -355 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -179 88 -145 104
rect -179 -104 -145 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 145 88 179 104
rect 145 -104 179 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 355 88 389 104
rect 355 -104 389 -88
rect 451 88 485 104
rect 451 -104 485 -88
rect -453 -181 -437 -147
rect -403 -181 -387 -147
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect 387 -181 403 -147
rect 437 -181 453 -147
rect -599 -249 -565 -187
rect 565 -249 599 -187
rect -599 -283 -503 -249
rect 503 -283 599 -249
<< viali >>
rect -227 147 -193 181
rect 193 147 227 181
rect -485 -88 -451 88
rect -389 -88 -355 88
rect -275 -88 -241 88
rect -179 -88 -145 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 145 -88 179 88
rect 241 -88 275 88
rect 355 -88 389 88
rect 451 -88 485 88
rect -437 -181 -403 -147
rect -17 -181 17 -147
rect 403 -181 437 -147
<< metal1 >>
rect -239 181 -181 187
rect -239 147 -227 181
rect -193 147 -181 181
rect -239 141 -181 147
rect 181 181 239 187
rect 181 147 193 181
rect 227 147 239 181
rect 181 141 239 147
rect -491 88 -445 100
rect -491 -88 -485 88
rect -451 -88 -445 88
rect -491 -100 -445 -88
rect -395 88 -349 100
rect -395 -88 -389 88
rect -355 -88 -349 88
rect -395 -100 -349 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -185 88 -139 100
rect -185 -88 -179 88
rect -145 -88 -139 88
rect -185 -100 -139 -88
rect -71 88 -25 100
rect -71 -88 -65 88
rect -31 -88 -25 88
rect -71 -100 -25 -88
rect 25 88 71 100
rect 25 -88 31 88
rect 65 -88 71 88
rect 25 -100 71 -88
rect 139 88 185 100
rect 139 -88 145 88
rect 179 -88 185 88
rect 139 -100 185 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 349 88 395 100
rect 349 -88 355 88
rect 389 -88 395 88
rect 349 -100 395 -88
rect 445 88 491 100
rect 445 -88 451 88
rect 485 -88 491 88
rect 445 -100 491 -88
rect -449 -147 -391 -141
rect -449 -181 -437 -147
rect -403 -181 -391 -147
rect -449 -187 -391 -181
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
rect 391 -147 449 -141
rect 391 -181 403 -147
rect 437 -181 449 -147
rect 391 -187 449 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -582 -266 582 266
string parameters w 1 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
