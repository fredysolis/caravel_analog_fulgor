**.subckt div_by_5 vdd vss CLK CLK_5 nCLK nQ2 Q1 Q0 nQ0 Q1_shift
*.iopin vdd
*.iopin vss
*.ipin CLK
*.opin CLK_5
*.ipin nCLK
*.iopin nQ2
*.iopin Q1
*.iopin Q0
*.iopin nQ0
*.iopin Q1_shift
x8 Q1 Q0 vss vss vdd vdd D2 sky130_fd_sc_hs__and2_1
x9 Q1 Q0 vss vss vdd vdd D1 sky130_fd_sc_hs__xor2_1
x10 nQ2 nQ0 vss vss vdd vdd D0 sky130_fd_sc_hs__and2_1
x12 Q1 Q1_shift vss vss vdd vdd CLK_5 sky130_fd_sc_hs__or2_1
x1 vdd Q2 nQ2 vss D2 CLK nCLK DFlipFlop
x2 vdd Q1 nQ1 vss D1 CLK nCLK DFlipFlop
x3 vdd Q0 nQ0 vss D0 CLK nCLK DFlipFlop
x4 vdd Q1_shift nQ1_shift vss Q1 nCLK CLK DFlipFlop
**.ends

* expanding   symbol:  DFlipFlop.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/DFlipFlop.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/DFlipFlop.sch
.subckt DFlipFlop  vdd Q nQ vss D CLK nCLK
*.iopin vdd
*.iopin vss
*.opin Q
*.opin nQ
*.ipin D
*.ipin CLK
*.ipin nCLK
x1 vdd D_d D nD_d vss clock_inverter
x2 vdd nA A D_d nD_d CLK vss latch_diff
x3 vdd nQ Q A nA nCLK vss latch_diff
.ends


* expanding   symbol:  clock_inverter.sym # of pins=5
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/clock_inverter.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/clock_inverter.sch
.subckt clock_inverter  vdd CLK_d CLK nCLK_d vss
*.ipin CLK
*.iopin vdd
*.iopin vss
*.opin nCLK_d
*.opin CLK_d
x5 vdd nCLK_d net1 vss trans_gate
x1 vdd CLK_d net2 vss inverter_cp_x1
x2 vdd net2 CLK vss inverter_cp_x1
x3 vdd net1 CLK vss inverter_cp_x1
.ends


* expanding   symbol:  latch_diff.sym # of pins=7
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/latch_diff.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/latch_diff.sch
.subckt latch_diff  vdd nQ Q D nD CLK vss
*.iopin vdd
*.iopin vss
*.ipin D
*.opin nQ
*.ipin CLK
*.ipin nD
*.opin Q
XM3 net1 CLK vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM4 nQ Q vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM5 Q nQ vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM1 nQ D net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 Q nD net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:  trans_gate.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/trans_gate.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/trans_gate.sch
.subckt trans_gate  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out vss in vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM1 out vdd in vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
.ends


* expanding   symbol:  inverter_cp_x1.sym # of pins=4
* sym_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_cp_x1.sym
* sch_path: /home/dhernando/caravel_analog_fulgor/xschem/inverter_cp_x1.sch
.subckt inverter_cp_x1  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
.ends

** flattened .save nodes
.end
