magic
tech sky130A
magscale 1 2
timestamp 1624402156
<< nwell >>
rect 19730 11269 20704 12071
rect 19753 11233 20704 11269
<< pwell >>
rect 14821 9774 17989 9782
rect 14905 9704 17989 9774
rect 14749 9518 14880 9540
rect 16610 9529 17989 9704
rect 16610 9518 17871 9529
rect 14749 9408 17871 9518
rect 14749 9262 17989 9408
<< ndiff >>
rect 19945 12469 20007 12481
rect 19945 12293 19957 12469
rect 19991 12293 20007 12469
rect 19945 12281 20007 12293
rect 20037 12469 20103 12481
rect 20037 12293 20053 12469
rect 20087 12293 20103 12469
rect 20037 12281 20103 12293
rect 20133 12469 20199 12481
rect 20133 12293 20149 12469
rect 20183 12293 20199 12469
rect 20133 12281 20199 12293
rect 20229 12469 20295 12481
rect 20229 12293 20245 12469
rect 20279 12293 20295 12469
rect 20229 12281 20295 12293
rect 20325 12469 20391 12481
rect 20325 12293 20341 12469
rect 20375 12293 20391 12469
rect 20325 12281 20391 12293
rect 20421 12469 20483 12481
rect 20421 12293 20437 12469
rect 20471 12293 20483 12469
rect 20421 12281 20483 12293
<< pdiff >>
rect 19868 11840 19926 11852
rect 19868 11464 19880 11840
rect 19914 11464 19926 11840
rect 19868 11452 19926 11464
rect 19996 11840 20054 11852
rect 19996 11464 20008 11840
rect 20042 11464 20054 11840
rect 19996 11452 20054 11464
rect 20124 11840 20182 11852
rect 20124 11464 20136 11840
rect 20170 11464 20182 11840
rect 20124 11452 20182 11464
rect 20252 11840 20310 11852
rect 20252 11464 20264 11840
rect 20298 11464 20310 11840
rect 20252 11452 20310 11464
rect 20380 11840 20438 11852
rect 20380 11464 20392 11840
rect 20426 11464 20438 11840
rect 20380 11452 20438 11464
rect 20508 11840 20566 11852
rect 20508 11464 20520 11840
rect 20554 11464 20566 11840
rect 20508 11452 20566 11464
<< ndiffc >>
rect 19957 12293 19991 12469
rect 20053 12293 20087 12469
rect 20149 12293 20183 12469
rect 20245 12293 20279 12469
rect 20341 12293 20375 12469
rect 20437 12293 20471 12469
<< pdiffc >>
rect 19880 11464 19914 11840
rect 20008 11464 20042 11840
rect 20136 11464 20170 11840
rect 20264 11464 20298 11840
rect 20392 11464 20426 11840
rect 20520 11464 20554 11840
<< locali >>
rect 19957 12469 19991 12485
rect 19957 12277 19991 12293
rect 20053 12469 20087 12485
rect 20053 12277 20087 12293
rect 20149 12469 20183 12485
rect 20149 12277 20183 12293
rect 20245 12469 20279 12485
rect 20245 12277 20279 12293
rect 20341 12469 20375 12485
rect 20341 12277 20375 12293
rect 20437 12469 20471 12485
rect 20437 12277 20471 12293
rect 19880 11840 19914 11856
rect 19880 11448 19914 11464
rect 20008 11840 20042 11856
rect 20008 11448 20042 11464
rect 20136 11840 20170 11856
rect 20136 11448 20170 11464
rect 20264 11840 20298 11856
rect 20264 11448 20298 11464
rect 20392 11840 20426 11856
rect 20392 11448 20426 11464
rect 20520 11840 20554 11856
rect 20520 11448 20554 11464
<< viali >>
rect 19920 12727 20470 12761
rect 19843 12621 20585 12655
rect 19957 12293 19991 12469
rect 20053 12293 20087 12469
rect 20149 12293 20183 12469
rect 20245 12293 20279 12469
rect 20341 12293 20375 12469
rect 20437 12293 20471 12469
rect 19880 11464 19914 11840
rect 20008 11464 20042 11840
rect 20136 11464 20170 11840
rect 20264 11464 20298 11840
rect 20392 11464 20426 11840
rect 20520 11464 20554 11840
rect 19766 11269 20668 11303
rect 19766 11163 20668 11197
rect 19843 9811 20585 9845
rect 19920 9705 20470 9739
<< metal1 >>
rect 14820 14616 18723 14756
rect 17273 13693 17300 13722
rect 14788 12514 17954 12991
rect 18583 12761 18723 14616
rect 20067 13133 20325 13283
rect 20028 12767 20074 12958
rect 20104 12901 20114 13101
rect 20180 12901 20190 13101
rect 20220 12767 20266 12963
rect 20296 12901 20306 13101
rect 20372 12901 20382 13101
rect 19908 12761 20482 12767
rect 18583 12727 19920 12761
rect 20470 12727 20585 12761
rect 18583 12661 20585 12727
rect 18583 12655 20597 12661
rect 18583 12621 19843 12655
rect 20585 12621 20597 12655
rect 19831 12615 20597 12621
rect 19099 12513 19105 12569
rect 19164 12513 20439 12569
rect 19951 12469 19997 12481
rect 19951 12293 19957 12469
rect 19991 12293 19997 12469
rect 19951 12141 19997 12293
rect 20027 12281 20037 12481
rect 20103 12281 20113 12481
rect 20143 12469 20189 12481
rect 20143 12293 20149 12469
rect 20183 12293 20189 12469
rect 20143 12141 20189 12293
rect 20219 12281 20229 12481
rect 20295 12281 20305 12481
rect 20335 12469 20381 12481
rect 20335 12293 20341 12469
rect 20375 12293 20381 12469
rect 20335 12141 20381 12293
rect 20411 12281 20421 12481
rect 20487 12281 20497 12481
rect 19273 12001 19283 12141
rect 19485 12001 20487 12141
rect 19874 11840 19920 12001
rect 19874 11464 19880 11840
rect 19914 11464 19920 11840
rect 19874 11452 19920 11464
rect 19986 11452 19996 11852
rect 20054 11452 20064 11852
rect 20130 11840 20176 12001
rect 20130 11464 20136 11840
rect 20170 11464 20176 11840
rect 20130 11452 20176 11464
rect 20242 11452 20252 11852
rect 20310 11452 20320 11852
rect 20386 11840 20432 12001
rect 20386 11464 20392 11840
rect 20426 11464 20432 11840
rect 20386 11452 20432 11464
rect 20498 11452 20508 11852
rect 20566 11452 20576 11852
rect 19605 11355 20508 11411
rect 19605 11261 19661 11355
rect 18246 11205 19661 11261
rect 19605 11111 19661 11205
rect 19754 11303 20680 11309
rect 19754 11269 19766 11303
rect 20668 11269 20680 11303
rect 20760 11269 20770 11290
rect 19754 11197 20770 11269
rect 19754 11163 19766 11197
rect 20668 11163 20680 11197
rect 20760 11180 20770 11197
rect 20864 11180 20874 11290
rect 19754 11157 20680 11163
rect 19605 11055 20508 11111
rect 19874 10465 19920 10793
rect 19986 10614 19996 11014
rect 20054 10614 20064 11014
rect 20130 10465 20176 10794
rect 20242 10614 20252 11014
rect 20310 10614 20320 11014
rect 20386 10465 20432 10789
rect 20498 10614 20508 11014
rect 20566 10614 20576 11014
rect 19273 10325 19283 10465
rect 19485 10325 20487 10465
rect 19951 10145 19997 10325
rect 14821 9934 15053 10037
rect 14821 9833 15499 9934
rect 17913 9890 19023 10037
rect 20027 9985 20037 10185
rect 20103 9985 20113 10185
rect 20143 10128 20189 10325
rect 20219 9985 20229 10185
rect 20295 9985 20305 10185
rect 20335 10146 20381 10325
rect 20411 9985 20421 10185
rect 20487 9985 20497 10185
rect 19099 9897 19105 9953
rect 19164 9897 20439 9953
rect 17883 9845 19023 9890
rect 19831 9845 20597 9851
rect 16103 9839 16629 9842
rect 17883 9839 19843 9845
rect 16103 9833 19843 9839
rect 14821 9811 19843 9833
rect 20585 9811 20597 9845
rect 14821 9805 20597 9811
rect 14821 9739 20585 9805
rect 14821 9705 19920 9739
rect 20470 9705 20585 9739
rect 14821 9701 19023 9705
rect 14821 9540 15170 9701
rect 15431 9540 15944 9701
rect 16205 9678 19023 9701
rect 19908 9699 20482 9705
rect 16205 9540 16635 9678
rect 16685 9644 19023 9678
rect 14036 9492 14176 9540
rect 14598 9528 16635 9540
rect 17883 9544 19023 9644
rect 20028 9546 20074 9699
rect 17883 9529 18500 9544
rect 14598 9518 14930 9528
rect 16469 9526 16635 9528
rect 14598 9516 15499 9518
rect 14821 9504 14930 9516
rect 15037 9512 15499 9516
rect 18314 9409 18500 9529
rect 20104 9365 20114 9565
rect 20180 9365 20190 9565
rect 20220 9558 20266 9699
rect 20296 9365 20306 9565
rect 20372 9365 20382 9565
rect 20067 9230 20325 9333
rect 17987 9050 18611 9058
rect 17987 8951 18047 9050
rect 18271 8951 18611 9050
rect 19066 8957 19076 9013
rect 19135 8957 19145 9013
rect 17987 8944 18611 8951
rect 5835 8187 6293 8311
rect 17989 8065 19076 8451
<< via1 >>
rect 20114 12901 20180 13101
rect 20306 12901 20372 13101
rect 19105 12513 19164 12569
rect 20037 12469 20103 12481
rect 20037 12293 20053 12469
rect 20053 12293 20087 12469
rect 20087 12293 20103 12469
rect 20037 12281 20103 12293
rect 20229 12469 20295 12481
rect 20229 12293 20245 12469
rect 20245 12293 20279 12469
rect 20279 12293 20295 12469
rect 20229 12281 20295 12293
rect 20421 12469 20487 12481
rect 20421 12293 20437 12469
rect 20437 12293 20471 12469
rect 20471 12293 20487 12469
rect 20421 12281 20487 12293
rect 19283 12001 19485 12141
rect 19996 11840 20054 11852
rect 19996 11464 20008 11840
rect 20008 11464 20042 11840
rect 20042 11464 20054 11840
rect 19996 11452 20054 11464
rect 20252 11840 20310 11852
rect 20252 11464 20264 11840
rect 20264 11464 20298 11840
rect 20298 11464 20310 11840
rect 20252 11452 20310 11464
rect 20508 11840 20566 11852
rect 20508 11464 20520 11840
rect 20520 11464 20554 11840
rect 20554 11464 20566 11840
rect 20508 11452 20566 11464
rect 20770 11180 20864 11290
rect 19996 10614 20054 11014
rect 20252 10614 20310 11014
rect 20508 10614 20566 11014
rect 19283 10325 19485 10465
rect 20037 9985 20103 10185
rect 20229 9985 20295 10185
rect 20421 9985 20487 10185
rect 19105 9897 19164 9953
rect 20114 9365 20180 9565
rect 20306 9365 20372 9565
rect 18047 8951 18271 9050
rect 19076 8957 19135 9013
<< metal2 >>
rect 14862 14658 14947 14708
rect 16088 13664 16201 13674
rect 16088 13529 16201 13539
rect 20114 13101 20180 13111
rect 20306 13101 20372 13111
rect 14788 12514 17954 12991
rect 20180 12901 20306 13101
rect 20372 12901 21067 13101
rect 20114 12891 20180 12901
rect 20306 12891 20372 12901
rect 19105 12569 19164 12579
rect 19105 12503 19164 12513
rect 15312 12422 15498 12432
rect 15312 12317 15498 12327
rect 14231 11343 14357 11411
rect 14231 11055 14357 11123
rect 6250 9575 6284 9607
rect 15061 9475 15095 9507
rect 18047 9050 18286 10381
rect 19109 9963 19160 12503
rect 20037 12481 20103 12491
rect 20229 12481 20295 12491
rect 20421 12481 20487 12491
rect 20867 12481 21067 12901
rect 20103 12281 20229 12481
rect 20295 12281 20421 12481
rect 20487 12281 21067 12481
rect 20037 12271 20103 12281
rect 20229 12271 20295 12281
rect 20421 12271 20487 12281
rect 19283 12141 19485 12151
rect 19283 11991 19485 12001
rect 19996 11852 20054 11862
rect 20252 11852 20310 11862
rect 20054 11568 20252 11768
rect 19996 11442 20054 11452
rect 20508 11852 20566 11862
rect 20310 11568 20508 11768
rect 20252 11442 20310 11452
rect 20867 11768 21067 12281
rect 20566 11568 21067 11768
rect 20508 11442 20566 11452
rect 20770 11293 20864 11300
rect 20770 11290 21302 11293
rect 20864 11182 21302 11290
rect 20770 11170 20864 11180
rect 19996 11014 20054 11024
rect 20252 11014 20310 11024
rect 20054 10698 20252 10898
rect 19996 10604 20054 10614
rect 20508 11014 20566 11024
rect 20310 10698 20508 10898
rect 20252 10604 20310 10614
rect 20566 10698 21067 10898
rect 20508 10604 20566 10614
rect 19283 10465 19485 10475
rect 19283 10315 19485 10325
rect 20037 10185 20103 10195
rect 20229 10185 20295 10195
rect 20421 10185 20487 10195
rect 20867 10185 21067 10698
rect 20103 9985 20229 10185
rect 20295 9985 20421 10185
rect 20487 9985 21067 10185
rect 20037 9975 20103 9985
rect 20229 9975 20295 9985
rect 20421 9975 20487 9985
rect 19105 9953 19164 9963
rect 19105 9887 19164 9897
rect 18271 8951 18286 9050
rect 19109 9023 19160 9887
rect 20114 9565 20180 9575
rect 20306 9565 20372 9575
rect 20867 9565 21067 9985
rect 20180 9365 20306 9565
rect 20372 9365 21067 9565
rect 20114 9355 20180 9365
rect 20210 9356 20276 9365
rect 20306 9355 20372 9365
rect 18047 8941 18286 8951
rect 19076 9013 19160 9023
rect 19135 8957 19160 9013
rect 19076 8947 19160 8957
<< via2 >>
rect 16088 13539 16201 13664
rect 15312 12327 15498 12422
rect 19283 12001 19485 12141
rect 19283 10325 19485 10465
<< metal3 >>
rect 16613 14055 16659 14110
rect 17217 14062 17263 14117
rect 18216 14056 18262 14111
rect 16082 13664 16211 13669
rect 16082 13539 16088 13664
rect 16201 13539 16211 13664
rect 16082 13534 16211 13539
rect 15303 12422 15508 12427
rect 15272 12327 15282 12422
rect 15498 12327 15508 12422
rect 15284 12317 15508 12327
rect 19273 12141 19495 12146
rect 19273 12001 19283 12141
rect 19485 12001 19495 12141
rect 19273 11996 19495 12001
rect 19273 10465 19495 10470
rect 19273 10325 19283 10465
rect 19485 10325 19495 10465
rect 19273 10320 19495 10325
rect 10019 9586 10053 9618
rect 5864 7650 5993 7651
rect 6199 7650 6259 7696
rect 5864 7590 6259 7650
rect 5864 7589 5993 7590
<< via3 >>
rect 16088 13539 16201 13664
rect 15282 12327 15312 12422
rect 15312 12327 15498 12422
rect 19283 12001 19485 12141
rect 19283 10325 19485 10465
<< metal4 >>
rect 15284 13665 16088 13669
rect 15284 13664 16202 13665
rect 15284 13539 16088 13664
rect 16201 13539 16202 13664
rect 15284 13538 16202 13539
rect 15284 13534 16088 13538
rect 15284 12423 15419 13534
rect 15281 12422 15499 12423
rect 15281 12327 15282 12422
rect 15498 12327 15499 12422
rect 15281 12326 15499 12327
rect 19282 12141 19486 12142
rect 19282 12001 19283 12141
rect 19485 12001 19486 12141
rect 19282 12000 19486 12001
rect 19283 11653 19485 12000
rect 18286 11451 19485 11653
rect 18084 10813 19485 11015
rect 19283 10466 19485 10813
rect 19282 10465 19486 10466
rect 19282 10325 19283 10465
rect 19485 10325 19486 10465
rect 19282 10324 19486 10325
rect 19283 10315 19485 10324
use inverter_min_x4  inverter_min_x4_0
timestamp 1624049879
transform 1 0 18411 0 -1 8928
box -53 -616 665 643
use res_amp_lin  res_amp_lin_0
timestamp 1624396448
transform 1 0 13177 0 1 11829
box 1054 -2058 5121 915
use delay_cell_buff  delay_cell_buff_0
timestamp 1624063007
transform 1 0 6173 0 1 7077
box -208 0 11816 2601
use sky130_fd_pr__nfet_01v8_lvt_72JNYZ  sky130_fd_pr__nfet_01v8_lvt_72JNYZ_0
timestamp 1624032293
transform 1 0 20195 0 -1 9465
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_lvt_595QY5  sky130_fd_pr__nfet_01v8_lvt_595QY5_0
timestamp 1624030292
transform 1 0 20214 0 1 10085
box -407 -310 407 310
use sky130_fd_pr__nfet_01v8_lvt_72JNYZ  sky130_fd_pr__nfet_01v8_lvt_72JNYZ_1
timestamp 1624032293
transform 1 0 20195 0 1 13001
box -311 -310 311 310
use sky130_fd_pr__pfet_01v8_lvt_4L9VGG  sky130_fd_pr__pfet_01v8_lvt_4L9VGG_0
timestamp 1624030292
transform 1 0 20217 0 1 10814
box -487 -419 487 419
use sky130_fd_pr__pfet_01v8_lvt_4L9VGG  sky130_fd_pr__pfet_01v8_lvt_4L9VGG_1
timestamp 1624030292
transform 1 0 20217 0 -1 11652
box -487 -419 487 419
use sky130_fd_pr__nfet_01v8_lvt_595QY5  sky130_fd_pr__nfet_01v8_lvt_595QY5_1
timestamp 1624030292
transform 1 0 20214 0 -1 12381
box -407 -310 407 310
use iref_ctrl_res_amp  iref_ctrl_res_amp_0
timestamp 1624113259
transform 1 0 15406 0 -1 14113
box -586 -686 2888 1369
<< labels >>
rlabel metal2 14231 11343 14357 11411 1 inn
rlabel metal2 14231 11055 14357 11123 1 inp
rlabel metal3 16613 14055 16659 14110 1 iref_reg0
rlabel metal3 17217 14062 17263 14117 1 iref_reg1
rlabel metal3 18216 14056 18262 14111 1 iref_reg2
rlabel metal1 17273 13693 17300 13722 1 iref
rlabel metal3 5878 7605 5911 7634 1 clk
rlabel metal2 6250 9575 6284 9607 1 delay_reg2
rlabel metal3 10019 9586 10053 9618 1 delay_reg1
rlabel metal2 15061 9475 15095 9507 1 delay_reg0
rlabel metal2 20931 12329 20986 12376 1 outp_cap
rlabel metal2 20931 10048 20986 10095 1 outn_cap
rlabel metal4 18370 10891 18425 10938 1 outn
rlabel metal4 18378 11537 18433 11584 1 outp
rlabel metal2 14898 14658 14947 14708 1 avss1p8
rlabel metal2 14841 12807 14890 12857 1 avdd1p8
rlabel metal1 20157 9238 20193 9270 1 rst
rlabel metal1 18156 8224 18193 8264 1 avdd1p8
rlabel metal1 20155 13197 20192 13237 1 rst
rlabel metal1 20715 11216 20746 11255 1 avdd1p8
<< end >>
