magic
tech sky130A
magscale 1 2
timestamp 1624653480
<< nwell >>
rect -64 618 579 637
rect -64 599 -17 618
rect -64 -47 -40 599
rect 568 -47 579 618
rect -64 -53 579 -47
<< pwell >>
rect -64 -725 579 -53
<< poly >>
rect 147 69 371 135
rect 279 30 371 69
rect 279 -34 301 30
rect 347 -34 371 30
rect 279 -53 371 -34
rect 145 -66 237 -53
rect 145 -130 168 -66
rect 214 -130 237 -66
rect 145 -171 237 -130
rect 145 -237 369 -171
<< polycont >>
rect 301 -34 347 30
rect 168 -130 214 -66
<< locali >>
rect 281 30 363 50
rect 281 -34 301 30
rect 347 -34 363 30
rect 151 -66 231 -48
rect 281 -57 363 -34
rect 151 -130 168 -66
rect 214 -130 231 -66
rect 151 -147 231 -130
<< viali >>
rect 79 565 437 599
rect 301 -34 347 30
rect 168 -130 214 -66
rect 79 -687 437 -653
<< metal1 >>
rect 67 599 449 605
rect 67 565 79 599
rect 437 565 449 599
rect 67 559 449 565
rect 45 490 329 508
rect -20 217 -10 490
rect 58 462 329 490
rect 58 404 137 462
rect 283 404 329 462
rect 58 217 97 404
rect 45 -171 97 217
rect 425 183 477 416
rect 187 120 233 178
rect 419 120 477 183
rect 187 74 477 120
rect 295 30 353 42
rect 285 -34 295 30
rect 353 -34 363 30
rect 295 -46 353 -34
rect 162 -66 220 -54
rect 152 -130 162 -66
rect 220 -130 230 -66
rect 162 -142 220 -130
rect 45 -217 329 -171
rect 45 -341 97 -217
rect 283 -263 329 -217
rect 419 -309 477 74
rect 45 -513 91 -341
rect 419 -343 465 -309
rect 425 -455 465 -343
rect 419 -501 465 -455
rect 187 -559 233 -513
rect 379 -559 465 -501
rect 187 -582 465 -559
rect 533 -582 543 -309
rect 187 -605 477 -582
rect 67 -653 449 -647
rect 67 -687 79 -653
rect 437 -687 449 -653
rect 67 -693 449 -687
<< via1 >>
rect -10 217 58 490
rect 295 -34 301 30
rect 301 -34 347 30
rect 347 -34 353 30
rect 162 -130 168 -66
rect 168 -130 214 -66
rect 214 -130 220 -66
rect 465 -582 533 -309
<< metal2 >>
rect -10 490 58 500
rect -10 207 58 217
rect 295 30 353 40
rect 295 -44 353 -34
rect 162 -66 220 -56
rect 162 -140 220 -130
rect 465 -309 533 -299
rect 465 -592 533 -582
<< via2 >>
rect -10 217 58 490
rect 465 -582 533 -309
<< metal3 >>
rect -20 490 68 495
rect -20 217 -10 490
rect 58 217 68 490
rect -20 212 68 217
rect 455 -309 543 -304
rect 455 -582 465 -309
rect 533 -582 543 -309
rect 455 -587 543 -582
use sky130_fd_pr__pfet_01v8_4798MH  sky130_fd_pr__pfet_01v8_4798MH_0
timestamp 1624062693
transform 1 0 258 0 1 291
box -311 -338 311 344
use sky130_fd_pr__nfet_01v8_BHR94T  sky130_fd_pr__nfet_01v8_BHR94T_0
timestamp 1624062693
transform 1 0 258 0 1 -388
box -311 -335 311 324
<< labels >>
rlabel metal1 67 -653 449 -647 1 vss
rlabel metal1 67 559 449 565 1 vdd
rlabel poly 279 -53 371 135 1 en_neg
rlabel poly 145 -237 237 -53 1 en_pos
rlabel metal1 419 -309 477 183 1 in
rlabel metal1 45 -341 97 217 1 out
<< end >>
