magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< metal1 >>
rect 0 1180 2872 1234
rect 0 652 210 718
rect 545 714 846 718
rect 545 662 791 714
rect 895 662 905 714
rect 1438 662 1448 714
rect 1552 662 1562 714
rect 545 652 846 662
rect 1979 652 2308 718
rect 1234 572 1244 624
rect 1348 572 1358 624
rect 256 497 266 549
rect 370 497 380 549
rect 896 472 906 524
rect 1010 472 1020 524
rect 1616 481 1626 533
rect 1730 481 1740 533
rect 2154 436 2220 557
rect 2680 481 2690 533
rect 2794 481 2804 533
rect 1949 380 1959 432
rect 2063 380 2073 432
rect 2149 332 2159 436
rect 2211 332 2221 436
rect 2154 329 2220 332
rect 0 70 2872 124
<< via1 >>
rect 791 662 895 714
rect 1448 662 1552 714
rect 1244 572 1348 624
rect 266 497 370 549
rect 906 472 1010 524
rect 1626 481 1730 533
rect 2690 481 2794 533
rect 1959 380 2063 432
rect 2159 332 2211 436
<< metal2 >>
rect 791 714 895 724
rect 1448 714 1552 724
rect 895 662 1448 714
rect 791 652 895 662
rect 1448 652 1552 662
rect 1244 624 1348 634
rect 266 572 1244 624
rect 1348 572 2872 624
rect 266 549 370 572
rect 1244 562 1348 572
rect 266 487 370 497
rect 906 524 1010 534
rect 906 462 1010 472
rect 1626 533 2794 543
rect 1730 491 2690 533
rect 1626 471 1730 481
rect 2690 471 2794 481
rect 931 432 983 462
rect 1959 432 2063 442
rect 931 380 1959 432
rect 1959 370 2063 380
rect 2159 436 2211 446
rect 2159 322 2211 332
use nor_pfd  nor_pfd_0
timestamp 1624049879
transform 1 0 235 0 1 -468
box -235 468 483 1772
use nor_pfd  nor_pfd_1
timestamp 1624049879
transform 1 0 953 0 1 -468
box -235 468 483 1772
use nor_pfd  nor_pfd_2
timestamp 1624049879
transform 1 0 1671 0 1 -468
box -235 468 483 1772
use nor_pfd  nor_pfd_3
timestamp 1624049879
transform 1 0 2389 0 1 -468
box -235 468 483 1772
<< labels >>
rlabel metal1 0 652 210 718 1 CLK
rlabel metal1 0 1180 2872 1234 1 vdd
rlabel metal1 0 70 2872 124 1 vss
rlabel metal2 2768 572 2872 624 1 Q
rlabel via1 2159 332 2211 436 1 Reset
<< end >>
