* NGSPICE file created from user_analog_prject_wrapper.ext - technology: sky130A


* Top level circuit user_analog_prject_wrapper

.end

