magic
tech sky130A
magscale 1 2
timestamp 1624397418
<< checkpaint >>
rect -4732 -4732 589003 708732
<< nwell >>
rect 14730 660108 64962 661110
rect 14730 660034 64841 660108
rect 82888 660083 133067 660649
rect 83408 660052 119178 660083
rect 14730 659150 14782 660034
rect 28401 659941 28758 659982
rect 83408 659846 112858 660052
rect 124441 660015 133067 660083
<< nsubdiff >>
rect 84063 660455 112263 660457
rect 23064 660357 28702 660375
rect 14777 660340 21696 660354
rect 14777 660170 14819 660340
rect 21653 660170 21696 660340
rect 14777 660157 21696 660170
rect 23064 660187 23112 660357
rect 28654 660187 28702 660357
rect 23064 660169 28702 660187
rect 28954 660354 34964 660367
rect 28954 660184 28984 660354
rect 34934 660184 34964 660354
rect 28954 660172 34964 660184
rect 35514 660346 63803 660369
rect 35514 660176 35565 660346
rect 63751 660176 63803 660346
rect 84063 660217 84104 660455
rect 112222 660217 112263 660455
rect 124754 660421 132564 660424
rect 119365 660387 124394 660416
rect 84063 660216 112263 660217
rect 35514 660153 63803 660176
rect 112659 660209 119108 660241
rect 112659 660107 112704 660209
rect 119062 660107 119108 660209
rect 119365 660217 119414 660387
rect 124344 660217 124394 660387
rect 119365 660188 124394 660217
rect 124754 660183 124800 660421
rect 132518 660183 132564 660421
rect 124754 660180 132564 660183
rect 112659 660076 119108 660107
<< nsubdiffcont >>
rect 14819 660170 21653 660340
rect 23112 660187 28654 660357
rect 28984 660184 34934 660354
rect 35565 660176 63751 660346
rect 84104 660217 112222 660455
rect 112704 660107 119062 660209
rect 119414 660217 124344 660387
rect 124800 660183 132518 660421
<< locali >>
rect 84071 660455 112255 660457
rect 23072 660361 28694 660375
rect 14785 660344 21688 660354
rect 14785 660340 14835 660344
rect 21637 660340 21688 660344
rect 14785 660170 14819 660340
rect 21653 660170 21688 660340
rect 14785 660166 14835 660170
rect 21637 660166 21688 660170
rect 23072 660183 23094 660361
rect 28672 660183 28694 660361
rect 23072 660169 28694 660183
rect 28962 660358 34956 660367
rect 28962 660354 28990 660358
rect 34928 660354 34956 660358
rect 28962 660184 28984 660354
rect 34934 660184 34956 660354
rect 28962 660180 28990 660184
rect 34928 660180 34956 660184
rect 28962 660172 34956 660180
rect 35522 660350 63795 660369
rect 35522 660172 35565 660350
rect 63751 660172 63795 660350
rect 84071 660217 84104 660455
rect 112222 660217 112255 660455
rect 124762 660421 132556 660424
rect 119373 660391 124386 660416
rect 84071 660216 112255 660217
rect 14785 660157 21688 660166
rect 35522 660153 63795 660172
rect 112667 660211 119100 660241
rect 112667 660105 112698 660211
rect 119068 660105 119100 660211
rect 119373 660213 119414 660391
rect 124344 660213 124386 660391
rect 119373 660188 124386 660213
rect 124762 660391 124800 660421
rect 132518 660391 132556 660421
rect 124762 660213 124790 660391
rect 132528 660213 132556 660391
rect 124762 660183 124800 660213
rect 132518 660183 132556 660213
rect 124762 660180 132556 660183
rect 112667 660076 119100 660105
<< viali >>
rect 14835 660340 21637 660344
rect 14835 660170 21637 660340
rect 14835 660166 21637 660170
rect 23094 660357 28672 660361
rect 23094 660187 23112 660357
rect 23112 660187 28654 660357
rect 28654 660187 28672 660357
rect 23094 660183 28672 660187
rect 28990 660354 34928 660358
rect 28990 660184 34928 660354
rect 28990 660180 34928 660184
rect 35565 660346 63751 660350
rect 35565 660176 63751 660346
rect 35565 660172 63751 660176
rect 84106 660247 112220 660425
rect 112698 660209 119068 660211
rect 112698 660107 112704 660209
rect 112704 660107 119062 660209
rect 119062 660107 119068 660209
rect 112698 660105 119068 660107
rect 119414 660387 124344 660391
rect 119414 660217 124344 660387
rect 119414 660213 124344 660217
rect 124790 660213 124800 660391
rect 124800 660213 132518 660391
rect 132518 660213 132528 660391
<< metal1 >>
rect 202956 688216 206559 688225
rect 202956 687844 202971 688216
rect 206543 687844 206559 688216
rect 202956 687835 206559 687844
rect 207113 688194 210605 688222
rect 207113 687822 207137 688194
rect 210581 687822 210605 688194
rect 207113 687795 210605 687822
rect 211166 688218 214658 688246
rect 211166 687846 211190 688218
rect 214634 687846 214658 688218
rect 227267 688245 230759 688273
rect 223050 688164 226874 688186
rect 223050 688060 223080 688164
rect 223016 687894 223080 688060
rect 211166 687819 214658 687846
rect 223050 687856 223080 687894
rect 226844 688060 226874 688164
rect 226844 687894 226915 688060
rect 226844 687856 226874 687894
rect 223050 687834 226874 687856
rect 227267 687873 227291 688245
rect 230735 687873 230759 688245
rect 227267 687846 230759 687873
rect 231320 688254 234812 688282
rect 231320 687882 231344 688254
rect 234788 687882 234812 688254
rect 231320 687855 234812 687882
rect 235302 688264 238794 688292
rect 235302 687892 235326 688264
rect 238770 687892 238794 688264
rect 235302 687865 238794 687892
rect 239323 688259 242815 688287
rect 239323 687887 239347 688259
rect 242791 687887 242815 688259
rect 239323 687860 242815 687887
rect 243362 688257 246854 688285
rect 243362 687885 243386 688257
rect 246830 687885 246854 688257
rect 243362 687858 246854 687885
rect 202763 685353 247155 685354
rect 202763 685045 202789 685353
rect 247129 685045 247155 685353
rect 202763 685044 247155 685045
rect 83775 660472 112339 660489
rect 83746 660453 112339 660472
rect 23004 660420 64063 660453
rect 23004 660397 23051 660420
rect 21700 660392 23051 660397
rect 14751 660356 23051 660392
rect 14751 660344 14859 660356
rect 14751 660166 14835 660344
rect 21637 660166 23051 660176
rect 14751 660112 23051 660166
rect 63999 660112 64063 660420
rect 14751 660070 64063 660112
rect 14751 660012 21718 660070
rect 23004 660030 64063 660070
rect 23037 660018 28912 660030
rect 83746 660017 83774 660453
rect 112306 660409 112339 660453
rect 119184 660429 133061 660493
rect 119184 660416 120283 660429
rect 112306 660408 112754 660409
rect 119106 660408 120283 660416
rect 112306 660391 120283 660408
rect 133007 660416 133061 660429
rect 112306 660328 119414 660391
rect 112306 660017 112671 660328
rect 119059 660213 119414 660328
rect 119059 660211 120283 660213
rect 119068 660121 120283 660211
rect 133007 660121 133067 660416
rect 119068 660105 133067 660121
rect 14751 659692 14783 660012
rect 83746 660010 112671 660017
rect 83746 659999 112334 660010
rect 112601 659956 112671 660010
rect 119059 660062 133067 660105
rect 119059 659956 119177 660062
rect 125643 660015 133067 660062
rect 112601 659944 119177 659956
rect 157073 659872 198016 659901
rect 157073 659500 157102 659872
rect 197986 659500 198016 659872
rect 157073 659472 198016 659500
rect 12990 659361 14703 659415
rect 12990 659117 13082 659361
rect 14606 659270 14703 659361
rect 133071 659297 133364 659303
rect 133071 659270 133095 659297
rect 14606 659204 14991 659270
rect 132917 659204 133095 659270
rect 14606 659117 14703 659204
rect 133071 659181 133095 659204
rect 133339 659181 133364 659297
rect 133071 659175 133364 659181
rect 12990 659070 14703 659117
rect 66160 659105 68592 659137
rect 66160 658984 66198 659105
rect 64423 658604 66198 658984
rect 63068 658320 66198 658604
rect 64423 657999 66198 658320
rect 66160 657901 66198 657999
rect 68554 658984 68592 659105
rect 68554 657999 68603 658984
rect 79846 658972 83253 658973
rect 79838 658952 83253 658972
rect 79838 658004 79868 658952
rect 82288 658604 83253 658952
rect 206575 658752 206868 658758
rect 206575 658728 206599 658752
rect 206248 658662 206599 658728
rect 206575 658636 206599 658662
rect 206843 658636 206868 658752
rect 206575 658630 206868 658636
rect 82288 658320 84035 658604
rect 149997 658524 156268 658555
rect 149987 658497 156268 658524
rect 82288 658004 83253 658320
rect 68554 657901 68592 657999
rect 79838 657988 83253 658004
rect 79838 657985 82318 657988
rect 66160 657870 68592 657901
rect 21150 657656 23650 657665
rect 21150 657540 21190 657656
rect 23610 657540 23650 657656
rect 124326 657657 126710 657669
rect 21150 657532 23650 657540
rect 64013 657266 64962 657593
rect 34969 657228 35070 657242
rect 34969 657176 34993 657228
rect 35045 657176 35070 657228
rect 34969 657163 35070 657176
rect 34989 656786 35045 657163
rect 34964 656759 35076 656786
rect 64135 656771 64962 657266
rect 64163 656761 64962 656771
rect 34964 656707 34994 656759
rect 35046 656707 35076 656759
rect 64457 656747 64962 656761
rect 82894 657275 83827 657583
rect 124326 657541 124340 657657
rect 126696 657541 126710 657657
rect 124326 657529 126710 657541
rect 149987 657421 150019 658497
rect 152311 658062 156268 658497
rect 152311 657778 157347 658062
rect 152311 657421 156268 657778
rect 149987 657395 156268 657421
rect 149997 657379 156268 657395
rect 34964 656680 35076 656707
rect 82894 656573 83702 657275
rect 112660 657227 112812 657243
rect 112660 657175 112678 657227
rect 112730 657175 112742 657227
rect 112794 657175 112812 657227
rect 112660 657160 112812 657175
rect 112685 656533 112741 657160
rect 197704 657121 199952 657125
rect 156207 656708 157418 657036
rect 197704 657005 197714 657121
rect 199942 657005 199952 657121
rect 197704 657001 199952 657005
rect 112626 656530 112807 656533
rect 112626 656350 112658 656530
rect 112774 656350 112807 656530
rect 112626 656348 112807 656350
rect 156207 656248 156786 656708
rect 186130 656688 186235 656702
rect 186130 656636 186156 656688
rect 186208 656636 186235 656688
rect 186130 656623 186235 656636
rect 186152 656414 186208 656623
rect 186119 656391 186251 656414
rect 186119 656339 186159 656391
rect 186211 656339 186251 656391
rect 186119 656316 186251 656339
rect 12125 655528 13406 655533
rect 12125 655200 14468 655528
rect 133382 655200 135242 655528
rect 12125 652870 13406 655200
rect 134093 653281 135239 655200
rect 207475 654986 208245 655013
rect 206694 654658 208245 654986
rect 12125 651670 15784 652870
rect 132088 652146 135239 653281
rect 207475 652403 208245 654658
rect 132558 652135 135239 652146
rect 12125 651669 15583 651670
rect 12125 651650 13406 651669
rect 205405 651403 208245 652403
rect 205405 651383 207885 651403
rect 124847 637259 125452 637281
rect 124847 637079 124867 637259
rect 125431 637079 125452 637259
rect 124847 637057 125452 637079
<< via1 >>
rect 202971 687844 206543 688216
rect 207137 687822 210581 688194
rect 211190 687846 214634 688218
rect 223080 687856 226844 688164
rect 227291 687873 230735 688245
rect 231344 687882 234788 688254
rect 235326 687892 238770 688264
rect 239347 687887 242791 688259
rect 243386 687885 246830 688257
rect 202789 685045 247129 685353
rect 23051 660361 63999 660420
rect 23051 660356 23094 660361
rect 14859 660344 23094 660356
rect 14859 660176 21637 660344
rect 21637 660183 23094 660344
rect 23094 660183 28672 660361
rect 28672 660358 63999 660361
rect 28672 660183 28990 660358
rect 21637 660180 28990 660183
rect 28990 660180 34928 660358
rect 34928 660350 63999 660358
rect 34928 660180 35565 660350
rect 21637 660176 35565 660180
rect 23051 660172 35565 660176
rect 35565 660172 63751 660350
rect 63751 660172 63999 660350
rect 23051 660112 63999 660172
rect 83774 660425 112306 660453
rect 83774 660247 84106 660425
rect 84106 660247 112220 660425
rect 112220 660247 112306 660425
rect 120283 660391 133007 660429
rect 83774 660017 112306 660247
rect 112671 660211 119059 660328
rect 120283 660213 124344 660391
rect 124344 660213 124790 660391
rect 124790 660213 132528 660391
rect 132528 660213 133007 660391
rect 112671 660105 112698 660211
rect 112698 660105 119059 660211
rect 120283 660121 133007 660213
rect 112671 659956 119059 660105
rect 157102 659500 197986 659872
rect 13082 659117 14606 659361
rect 133095 659181 133339 659297
rect 66198 657901 68554 659105
rect 79868 658004 82288 658952
rect 206599 658636 206843 658752
rect 21190 657540 23610 657656
rect 34993 657176 35045 657228
rect 34994 656707 35046 656759
rect 124340 657541 126696 657657
rect 150019 657421 152311 658497
rect 112678 657175 112730 657227
rect 112742 657175 112794 657227
rect 197714 657005 199942 657121
rect 112658 656350 112774 656530
rect 186156 656636 186208 656688
rect 186159 656339 186211 656391
rect 124867 637079 125431 637259
<< metal2 >>
rect 211169 688677 214642 688713
rect 207123 688597 210596 688633
rect 198295 688226 199269 688229
rect 202966 688226 206549 688235
rect 198295 688216 206549 688226
rect 198295 688212 202971 688216
rect 198295 687836 198314 688212
rect 199250 687844 202971 688212
rect 206543 687844 206549 688216
rect 199250 687836 206549 687844
rect 198295 687825 206549 687836
rect 207123 688194 207151 688597
rect 210567 688194 210596 688597
rect 198295 687820 199269 687825
rect 207123 687822 207137 688194
rect 210581 687822 210596 688194
rect 211169 688218 211197 688677
rect 214613 688256 214642 688677
rect 227277 688638 230750 688674
rect 214613 688218 214648 688256
rect 211169 687865 211190 688218
rect 207123 687821 207151 687822
rect 210567 687821 210596 687822
rect 207123 687785 210596 687821
rect 211176 687846 211190 687865
rect 214634 687846 214648 688218
rect 227277 688245 227305 688638
rect 230721 688245 230750 688638
rect 211176 687809 214648 687846
rect 223060 688164 226864 688196
rect 223060 687856 223080 688164
rect 226844 687856 226864 688164
rect 223060 687824 226864 687856
rect 227277 687873 227291 688245
rect 230735 687873 230750 688245
rect 227277 687862 227305 687873
rect 230721 687862 230750 687873
rect 227277 687826 230750 687862
rect 231330 688657 234803 688693
rect 231330 688254 231358 688657
rect 234774 688254 234803 688657
rect 231330 687882 231344 688254
rect 234788 687882 234803 688254
rect 231330 687881 231358 687882
rect 234774 687881 234803 687882
rect 231330 687845 234803 687881
rect 235312 688667 238785 688703
rect 235312 688264 235340 688667
rect 238756 688264 238785 688667
rect 235312 687892 235326 688264
rect 238770 687892 238785 688264
rect 235312 687891 235340 687892
rect 238756 687891 238785 687892
rect 235312 687855 238785 687891
rect 239333 688662 242806 688698
rect 239333 688259 239361 688662
rect 242777 688259 242806 688662
rect 239333 687887 239347 688259
rect 242791 687887 242806 688259
rect 239333 687886 239361 687887
rect 242777 687886 242806 687887
rect 239333 687850 242806 687886
rect 243372 688660 246845 688696
rect 243372 688257 243400 688660
rect 246816 688257 246845 688660
rect 243372 687885 243386 688257
rect 246830 687885 246845 688257
rect 243372 687884 243400 687885
rect 246816 687884 246845 687885
rect 243372 687848 246845 687884
rect 202773 685353 247145 685364
rect 202773 685045 202789 685353
rect 247129 685045 247145 685353
rect 202773 685034 202813 685045
rect 202780 684733 202813 685034
rect 247109 685034 247145 685045
rect 247109 684733 247142 685034
rect 202780 684701 247142 684733
rect 83765 660820 124085 660856
rect 23042 660647 64025 660667
rect 23042 660420 23065 660647
rect 23042 660398 23051 660420
rect 14834 660356 23051 660398
rect 14834 660176 14859 660356
rect 14834 660112 23051 660176
rect 14834 660111 23065 660112
rect 64001 660111 64025 660647
rect 83765 660482 83777 660820
rect 23042 660091 64025 660111
rect 83756 660453 83777 660482
rect 124073 660455 124085 660820
rect 157083 660495 197708 660512
rect 83756 660017 83774 660453
rect 124073 660429 133038 660455
rect 112306 660017 112671 660204
rect 83756 659999 112671 660017
rect 83756 659989 112324 659999
rect 112657 659956 112671 659999
rect 119059 660121 120283 660204
rect 133007 660121 133038 660429
rect 119059 660096 133038 660121
rect 119059 659999 120418 660096
rect 119059 659956 119074 659999
rect 112657 659943 119074 659956
rect 2509 659751 14155 659826
rect 2509 658735 2684 659751
rect 5060 659386 14155 659751
rect 133210 659530 140004 659630
rect 5060 659361 14624 659386
rect 5060 659117 13082 659361
rect 14606 659117 14624 659361
rect 133210 659313 137615 659530
rect 133081 659297 137615 659313
rect 133081 659181 133095 659297
rect 133339 659181 137615 659297
rect 133081 659165 137615 659181
rect 5060 659093 14624 659117
rect 66170 659131 68582 659147
rect 5060 658735 14155 659093
rect 2509 658656 14155 658735
rect 66170 657875 66188 659131
rect 68564 657875 68582 659131
rect 79848 658952 82308 658982
rect 79848 658946 79868 658952
rect 82288 658946 82308 658952
rect 79848 658010 79850 658946
rect 82306 658010 82308 658946
rect 133210 658914 137615 659165
rect 139911 658914 140004 659530
rect 157083 659479 157087 660495
rect 197703 659911 197708 660495
rect 197703 659872 198006 659911
rect 197986 659500 198006 659872
rect 197703 659479 198006 659500
rect 157083 659462 198006 659479
rect 133210 658850 140004 658914
rect 206714 659004 212383 659085
rect 206714 658768 209991 659004
rect 206585 658752 209991 658768
rect 206585 658636 206599 658752
rect 206843 658636 209991 658752
rect 206585 658620 209991 658636
rect 79848 658004 79868 658010
rect 82288 658004 82308 658010
rect 79848 657975 82308 658004
rect 149997 658507 152333 658534
rect 66170 657860 68582 657875
rect 21160 657679 23631 657700
rect 21160 657543 21167 657679
rect 23623 657675 23631 657679
rect 23623 657543 23640 657675
rect 21160 657540 21190 657543
rect 23610 657540 23640 657543
rect 21160 657522 23640 657540
rect 124336 657667 126700 657679
rect 124336 657657 124370 657667
rect 126666 657657 126700 657667
rect 124336 657541 124340 657657
rect 126696 657541 126700 657657
rect 124336 657531 124370 657541
rect 126666 657531 126700 657541
rect 124336 657519 126700 657531
rect 149997 657411 150017 658507
rect 152313 657411 152333 658507
rect 206714 658388 209991 658620
rect 212287 658388 212383 659004
rect 206714 658305 212383 658388
rect 149997 657385 152333 657411
rect 34979 657233 35060 657252
rect 32682 657228 35060 657233
rect 32682 657177 34993 657228
rect 34979 657176 34993 657177
rect 35045 657176 35060 657228
rect 34979 657153 35060 657176
rect 112670 657233 112802 657253
rect 112670 657227 115172 657233
rect 112670 657175 112678 657227
rect 112730 657175 112742 657227
rect 112794 657177 115172 657227
rect 112794 657175 112802 657177
rect 112670 657150 112802 657175
rect 197714 657121 199942 657135
rect 73065 657013 74069 657038
rect 73065 656798 73099 657013
rect 34974 656766 35066 656796
rect 35452 656766 73099 656798
rect 34974 656759 73099 656766
rect 34974 656707 34994 656759
rect 35046 656710 73099 656759
rect 35046 656707 35066 656710
rect 34974 656670 35066 656707
rect 35452 656678 73099 656710
rect 73065 656237 73099 656678
rect 74035 656488 74069 657013
rect 197714 656991 199942 657005
rect 186140 656691 186225 656712
rect 186140 656688 188420 656691
rect 186140 656636 186156 656688
rect 186208 656636 188420 656688
rect 186140 656635 188420 656636
rect 186140 656613 186225 656635
rect 112636 656530 112797 656543
rect 112636 656488 112658 656530
rect 74035 656363 112658 656488
rect 74035 656237 74069 656363
rect 112636 656350 112658 656363
rect 112774 656350 112797 656530
rect 112636 656338 112797 656350
rect 152623 656393 186037 656431
rect 186129 656393 186241 656424
rect 152623 656391 186241 656393
rect 152623 656376 186159 656391
rect 152623 656300 152664 656376
rect 73065 656212 74069 656237
rect 152633 656160 152664 656300
rect 153760 656339 186159 656376
rect 186211 656339 186241 656391
rect 153760 656337 186241 656339
rect 153760 656300 186037 656337
rect 186129 656306 186241 656337
rect 153760 656160 153791 656300
rect 152633 656124 153791 656160
rect 144160 637398 145498 637413
rect 144160 637369 144161 637398
rect 125227 637291 144161 637369
rect 124857 637259 144161 637291
rect 124857 637079 124867 637259
rect 125431 637079 144161 637259
rect 124857 637047 144161 637079
rect 125227 636972 144161 637047
rect 144160 636942 144161 636972
rect 145497 637369 145498 637398
rect 145497 636972 145544 637369
rect 145497 636942 145498 636972
rect 144160 636927 145498 636942
rect 368681 635496 368816 635526
rect 368681 635440 368720 635496
rect 368776 635440 368816 635496
rect 368681 635411 368816 635440
rect 368680 633658 368815 633688
rect 368680 633602 368719 633658
rect 368775 633602 368815 633658
rect 368680 633573 368815 633602
rect 152624 510668 153820 510686
rect 152624 510561 152634 510668
rect 1323 510535 152634 510561
rect 1323 510239 1376 510535
rect 2152 510508 152634 510535
rect 2152 510292 73033 510508
rect 74049 510292 152634 510508
rect 2152 510239 152634 510292
rect 1323 510212 152634 510239
rect 153810 510561 153820 510668
rect 153810 510212 153853 510561
rect 152624 510195 153820 510212
rect 1326 467314 145524 467339
rect 1326 467313 144193 467314
rect 1326 467017 1379 467313
rect 2155 467018 144193 467313
rect 145449 467018 145524 467314
rect 2155 467017 145524 467018
rect 1326 466990 145524 467017
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 198314 687836 199250 688212
rect 207151 688194 210567 688597
rect 207151 687822 210567 688194
rect 211197 688218 214613 688677
rect 211197 687901 214613 688218
rect 207151 687821 210567 687822
rect 227305 688245 230721 688638
rect 223094 687862 226830 688158
rect 227305 687873 230721 688245
rect 227305 687862 230721 687873
rect 231358 688254 234774 688657
rect 231358 687882 234774 688254
rect 231358 687881 234774 687882
rect 235340 688264 238756 688667
rect 235340 687892 238756 688264
rect 235340 687891 238756 687892
rect 239361 688259 242777 688662
rect 239361 687887 242777 688259
rect 239361 687886 242777 687887
rect 243400 688257 246816 688660
rect 243400 687885 246816 688257
rect 243400 687884 246816 687885
rect 202813 685045 247109 685269
rect 202813 684733 247109 685045
rect 23065 660420 64001 660647
rect 23065 660112 63999 660420
rect 63999 660112 64001 660420
rect 23065 660111 64001 660112
rect 83777 660453 124073 660820
rect 83777 660204 112306 660453
rect 112306 660429 124073 660453
rect 112306 660328 120283 660429
rect 112306 660204 112671 660328
rect 112671 660204 119059 660328
rect 119059 660204 120283 660328
rect 120283 660204 124073 660429
rect 2684 658735 5060 659751
rect 66188 659105 68564 659131
rect 66188 657901 66198 659105
rect 66198 657901 68554 659105
rect 68554 657901 68564 659105
rect 66188 657875 68564 657901
rect 79850 658010 79868 658946
rect 79868 658010 82288 658946
rect 82288 658010 82306 658946
rect 137615 658914 139911 659530
rect 157087 659872 197703 660495
rect 157087 659500 157102 659872
rect 157102 659500 197703 659872
rect 157087 659479 197703 659500
rect 21167 657656 23623 657679
rect 21167 657543 21190 657656
rect 21190 657543 23610 657656
rect 23610 657543 23623 657656
rect 124370 657657 126666 657667
rect 124370 657541 126666 657657
rect 124370 657531 126666 657541
rect 150017 658497 152313 658507
rect 150017 657421 150019 658497
rect 150019 657421 152311 658497
rect 152311 657421 152313 658497
rect 150017 657411 152313 657421
rect 209991 658388 212287 659004
rect 73099 656237 74035 657013
rect 197720 657035 197776 657091
rect 197800 657035 197856 657091
rect 197880 657035 197936 657091
rect 197960 657035 198016 657091
rect 198040 657035 198096 657091
rect 198120 657035 198176 657091
rect 198200 657035 198256 657091
rect 198280 657035 198336 657091
rect 198360 657035 198416 657091
rect 198440 657035 198496 657091
rect 198520 657035 198576 657091
rect 198600 657035 198656 657091
rect 198680 657035 198736 657091
rect 198760 657035 198816 657091
rect 198840 657035 198896 657091
rect 198920 657035 198976 657091
rect 199000 657035 199056 657091
rect 199080 657035 199136 657091
rect 199160 657035 199216 657091
rect 199240 657035 199296 657091
rect 199320 657035 199376 657091
rect 199400 657035 199456 657091
rect 199480 657035 199536 657091
rect 199560 657035 199616 657091
rect 199640 657035 199696 657091
rect 199720 657035 199776 657091
rect 199800 657035 199856 657091
rect 199880 657035 199936 657091
rect 152664 656160 153760 656376
rect 144161 636942 145497 637398
rect 368720 635440 368776 635496
rect 368719 633602 368775 633658
rect 1376 510239 2152 510535
rect 73033 510292 74049 510508
rect 152634 510212 153810 510668
rect 1379 467017 2155 467313
rect 144193 467018 145449 467314
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 704716 515394 704800
rect 520594 704716 525394 704800
rect 510296 704677 525583 704716
rect 17496 693341 19996 702300
rect 69842 699968 72342 702300
rect 69842 697468 82326 699968
rect 17498 693225 19996 693341
rect 17498 690841 17558 693225
rect 19942 690841 19996 693225
rect 17498 690746 19996 690841
rect 66130 693220 68630 693269
rect 66130 690836 66218 693220
rect 68522 690836 68630 693220
rect -800 683796 1700 685242
rect 21882 683875 22864 683906
rect -800 681296 5105 683796
rect 21882 681731 21901 683875
rect 22845 681731 22864 683875
rect 21882 681701 22864 681731
rect -800 680242 1700 681296
rect 2605 659751 5105 681296
rect 2605 658735 2684 659751
rect 5060 658735 5105 659751
rect -800 643842 1660 648642
rect -800 633842 1660 638642
rect 2605 611721 5105 658735
rect 21889 657695 22824 681701
rect 23032 661237 64027 661269
rect 23032 660133 23057 661237
rect 64001 660662 64027 661237
rect 23032 660111 23065 660133
rect 64001 660111 64035 660662
rect 23032 660096 64035 660111
rect 66130 659131 68630 690836
rect 66130 657875 66188 659131
rect 68564 657875 68630 659131
rect 79826 658946 82326 697468
rect 121407 699624 123907 702300
rect 121407 697124 152455 699624
rect 93805 695840 95820 695904
rect 93805 693936 93859 695840
rect 95763 693936 95820 695840
rect 93805 683877 95820 693936
rect 124995 692284 125965 692310
rect 124995 692109 125008 692284
rect 93805 681853 93870 683877
rect 93833 681813 93870 681853
rect 95694 681853 95820 683877
rect 124989 690380 125008 692109
rect 125952 690380 125965 692284
rect 124989 690355 125965 690380
rect 95694 681813 95731 681853
rect 93833 681797 95731 681813
rect 83755 661465 124081 661487
rect 83755 660201 83766 661465
rect 124070 660851 124081 661465
rect 124070 660820 124095 660851
rect 124073 660204 124095 660820
rect 124070 660201 124095 660204
rect 83755 660174 124095 660201
rect 79826 658010 79850 658946
rect 82306 658010 82326 658946
rect 79826 657959 82326 658010
rect 21150 657679 23641 657695
rect 21150 657543 21167 657679
rect 23623 657543 23641 657679
rect 66130 657635 68630 657875
rect 124989 657674 125924 690355
rect 137480 659530 139980 659593
rect 137480 658914 137615 659530
rect 139911 658914 139980 659530
rect 124326 657667 126710 657674
rect 21150 657527 23641 657543
rect 124326 657531 124370 657667
rect 126666 657531 126710 657667
rect 124326 657524 126710 657531
rect 72999 657013 74122 657160
rect 72999 656237 73099 657013
rect 74035 656237 74122 657013
rect 14417 624595 64654 624619
rect 14417 621651 14463 624595
rect 64607 621651 64654 624595
rect 14417 621627 64654 621651
rect 2605 607134 2674 611721
rect 2636 607097 2674 607134
rect 4978 607134 5105 611721
rect 4978 607097 5017 607134
rect 2636 607093 5017 607097
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect -800 511530 480 511642
rect 1348 510535 2181 510543
rect 1348 510460 1376 510535
rect -800 510348 1376 510460
rect 1292 510340 1376 510348
rect 1348 510239 1376 510340
rect 2152 510239 2181 510535
rect 1348 510231 2181 510239
rect 72999 510508 74122 656237
rect 83142 624590 133420 624630
rect 83142 622046 83169 624590
rect 133393 622046 133420 624590
rect 83142 622007 133420 622046
rect 137480 611815 139980 658914
rect 149955 658507 152455 697124
rect 166763 695391 169263 702300
rect 177015 695391 179515 702300
rect 218640 697297 221140 702300
rect 166762 692889 179515 695391
rect 211648 695751 214101 695778
rect 211648 694007 211682 695751
rect 214066 695500 214101 695751
rect 214066 694007 214151 695500
rect 218640 694913 218739 697297
rect 221043 694913 221140 697297
rect 218640 694879 221140 694913
rect 223860 697326 226360 697368
rect 223860 694942 223943 697326
rect 226247 694942 226360 697326
rect 211648 693981 214151 694007
rect 171983 684070 174483 692889
rect 207536 692333 210036 692388
rect 207536 690349 207618 692333
rect 209922 690349 210036 692333
rect 207536 688628 210036 690349
rect 211651 688708 214151 693981
rect 211159 688677 214652 688708
rect 207113 688597 210606 688628
rect 198292 688224 199274 688239
rect 198285 688212 199279 688224
rect 198285 687836 198314 688212
rect 199250 687836 199279 688212
rect 198285 687825 199279 687836
rect 171983 681570 192882 684070
rect 190382 667305 192882 681570
rect 190367 667282 192884 667305
rect 190367 664818 190393 667282
rect 192857 664818 192884 667282
rect 190367 664796 192884 664818
rect 157073 660499 197718 660507
rect 157073 659475 157083 660499
rect 197707 659475 197718 660499
rect 157073 659467 197718 659475
rect 149955 657411 150017 658507
rect 152313 657411 152455 658507
rect 149955 657301 152455 657411
rect 198292 657130 199274 687825
rect 207113 687821 207151 688597
rect 210567 687821 210606 688597
rect 211159 687901 211197 688677
rect 214613 687901 214652 688677
rect 223860 688191 226360 694942
rect 228892 697340 231392 702300
rect 242722 702116 245242 702134
rect 242722 699652 242750 702116
rect 245214 702114 245242 702116
rect 245214 699652 315546 702114
rect 242722 699634 315546 699652
rect 243372 699614 315546 699634
rect 228892 694956 228987 697340
rect 231291 694956 231392 697340
rect 228892 694833 231392 694956
rect 232116 696758 311894 699258
rect 232116 688688 234616 696758
rect 235915 693974 307678 696474
rect 235915 688698 238415 693974
rect 239738 691142 303725 693642
rect 227267 688661 230760 688669
rect 211159 687870 214652 687901
rect 223050 688158 226874 688191
rect 223050 687862 223094 688158
rect 226830 687862 226874 688158
rect 223050 687829 226874 687862
rect 227267 688117 227301 688661
rect 230725 688117 230760 688661
rect 227267 687862 227305 688117
rect 230721 687862 230760 688117
rect 227267 687831 230760 687862
rect 231320 688657 234813 688688
rect 231320 687881 231358 688657
rect 234774 687881 234813 688657
rect 231320 687850 234813 687881
rect 235302 688667 238795 688698
rect 239738 688693 242238 691142
rect 235302 687891 235340 688667
rect 238756 687891 238795 688667
rect 235302 687860 238795 687891
rect 239323 688662 242816 688693
rect 239323 687886 239361 688662
rect 242777 687886 242816 688662
rect 239323 687855 242816 687886
rect 243362 688660 299390 690785
rect 243362 687884 243400 688660
rect 246816 688285 299390 688660
rect 246816 687884 246855 688285
rect 243362 687853 246855 687884
rect 207113 687790 210606 687821
rect 202770 685278 247152 685296
rect 202770 684706 202809 685278
rect 247113 684734 247152 685278
rect 247109 684733 247152 684734
rect 202795 684094 202809 684706
rect 247033 684706 247152 684733
rect 247033 684094 247119 684706
rect 202795 684082 247119 684094
rect 209899 659004 212399 659121
rect 209899 658388 209991 659004
rect 212287 658388 212399 659004
rect 197704 657091 199952 657130
rect 197704 657035 197720 657091
rect 197776 657035 197800 657091
rect 197856 657035 197880 657091
rect 197936 657035 197960 657091
rect 198016 657035 198040 657091
rect 198096 657035 198120 657091
rect 198176 657035 198200 657091
rect 198256 657035 198280 657091
rect 198336 657035 198360 657091
rect 198416 657035 198440 657091
rect 198496 657035 198520 657091
rect 198576 657035 198600 657091
rect 198656 657035 198680 657091
rect 198736 657035 198760 657091
rect 198816 657035 198840 657091
rect 198896 657035 198920 657091
rect 198976 657035 199000 657091
rect 199056 657035 199080 657091
rect 199136 657035 199160 657091
rect 199216 657035 199240 657091
rect 199296 657035 199320 657091
rect 199376 657035 199400 657091
rect 199456 657035 199480 657091
rect 199536 657035 199560 657091
rect 199616 657035 199640 657091
rect 199696 657035 199720 657091
rect 199776 657035 199800 657091
rect 199856 657035 199880 657091
rect 199936 657035 199952 657091
rect 197704 656996 199952 657035
rect 152609 656376 153837 656431
rect 152609 656160 152664 656376
rect 153760 656160 153837 656376
rect 137480 607191 137770 611815
rect 139754 607191 139980 611815
rect 137480 607076 139980 607191
rect 144145 637398 145521 637418
rect 144145 636942 144161 637398
rect 145497 636942 145521 637398
rect 72999 510292 73033 510508
rect 74049 510292 74122 510508
rect 72999 510192 74122 510292
rect -800 509166 480 509278
rect -800 507984 490 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect 1351 467313 2184 467321
rect -800 467230 480 467238
rect 1351 467230 1379 467313
rect -800 467126 1379 467230
rect 304 467118 1379 467126
rect 1351 467017 1379 467118
rect 2155 467017 2184 467313
rect 1351 467009 2184 467017
rect 144145 467314 145521 636942
rect 152609 510668 153837 656160
rect 156490 624090 206846 624128
rect 156490 620746 156516 624090
rect 206820 620746 206846 624090
rect 156490 620709 206846 620746
rect 209899 611719 212399 658388
rect 296890 658340 299390 688285
rect 301225 661655 303725 691142
rect 305178 664670 307678 693974
rect 309394 668158 311894 696758
rect 313046 671728 315546 699614
rect 320335 695123 322835 702300
rect 330587 695123 333087 702300
rect 414564 696421 417064 702300
rect 466720 696421 469220 702300
rect 510296 701813 510307 704677
rect 510296 701790 510467 701813
rect 510456 697733 510467 701790
rect 525571 697733 525583 704677
rect 566594 702300 571594 704800
rect 567875 698736 570375 702300
rect 510456 697694 525583 697733
rect 567865 698718 570385 698736
rect 567865 696734 567893 698718
rect 570357 696734 570385 698718
rect 567865 696717 570385 696734
rect 320334 692621 333087 695123
rect 414554 696403 417074 696421
rect 414554 693939 414582 696403
rect 417046 693939 417074 696403
rect 414554 693921 417074 693939
rect 466710 696403 469230 696421
rect 466710 693939 466738 696403
rect 469202 693939 469230 696403
rect 466710 693921 469230 693939
rect 313036 671710 315556 671728
rect 313036 669246 313064 671710
rect 315528 669246 315556 671710
rect 313036 669228 315556 669246
rect 309384 668140 311904 668158
rect 309384 665676 309412 668140
rect 311876 665676 311904 668140
rect 309384 665658 311904 665676
rect 305168 664652 307688 664670
rect 305168 662188 305196 664652
rect 307660 662188 307688 664652
rect 305168 662170 307688 662188
rect 301215 661637 303735 661655
rect 301215 659173 301243 661637
rect 303707 659173 303735 661637
rect 301215 659155 303735 659173
rect 296880 658322 299400 658340
rect 296880 655858 296908 658322
rect 299372 655858 299400 658322
rect 296880 655840 299400 655858
rect 325555 650863 328055 692621
rect 582300 681668 584800 682984
rect 576277 681650 584800 681668
rect 576277 679186 576304 681650
rect 578288 679186 584800 681650
rect 576277 679168 584800 679186
rect 582300 677984 584800 679168
rect 373465 671710 374835 671728
rect 373465 669246 373478 671710
rect 374822 669246 374835 671710
rect 373465 669228 374835 669246
rect 371778 668140 373148 668158
rect 371778 665676 371791 668140
rect 373135 665676 373148 668140
rect 371778 665658 373148 665676
rect 369963 664652 371333 664670
rect 369963 662188 369976 664652
rect 371320 662188 371333 664652
rect 369963 662170 371333 662188
rect 368199 661655 369549 661704
rect 368189 661637 369559 661655
rect 368189 659173 368202 661637
rect 369546 659173 369559 661637
rect 368189 659155 369559 659173
rect 366150 658322 367520 658340
rect 366150 655858 366163 658322
rect 367507 655858 367520 658322
rect 366150 655840 367520 655858
rect 325545 650845 328065 650863
rect 325545 648381 325573 650845
rect 328037 648381 328065 650845
rect 325545 648363 328065 648381
rect 325555 648358 328055 648363
rect 366160 642905 367510 655840
rect 368199 642905 369549 659155
rect 369973 642905 371323 662170
rect 371788 642905 373138 665658
rect 373475 642905 374825 669228
rect 367006 642208 367202 642905
rect 360862 642012 367202 642208
rect 347630 637114 348966 637147
rect 347630 636730 347669 637114
rect 348053 636730 348966 637114
rect 360862 636883 361058 642012
rect 368630 641752 368826 642905
rect 368630 641556 370520 641752
rect 347630 636697 348966 636730
rect 368671 635496 368826 635521
rect 368671 635440 368720 635496
rect 368776 635440 368826 635496
rect 368671 635418 368826 635440
rect 368652 635049 368848 635418
rect 370324 635049 370520 641556
rect 368652 634853 370520 635049
rect 370918 634243 371114 642905
rect 372372 642103 372568 642905
rect 371439 641907 372568 642103
rect 371439 637006 371635 641907
rect 374402 641653 374598 642905
rect 371879 641457 374598 641653
rect 368651 634047 371114 634243
rect 368651 633658 368847 634047
rect 368651 633602 368719 633658
rect 368775 633602 368847 633658
rect 368651 633588 368847 633602
rect 368670 633578 368825 633588
rect 371879 632836 372075 641457
rect 582340 639784 584800 644584
rect 371440 632640 372075 632836
rect 371440 632181 371636 632640
rect 352226 630274 352712 630281
rect 352226 630050 352237 630274
rect 352701 630050 352712 630274
rect 358816 630277 359302 630284
rect 352226 613751 352712 630050
rect 356365 630255 356851 630262
rect 356365 630031 356376 630255
rect 356840 630031 356851 630255
rect 356365 615037 356851 630031
rect 358816 630053 358827 630277
rect 359291 630053 359302 630277
rect 358816 616322 359302 630053
rect 582340 629784 584800 634584
rect 361089 628732 361575 628785
rect 360254 628619 360672 628648
rect 360218 628609 360704 628619
rect 360218 628385 360271 628609
rect 360655 628385 360704 628609
rect 360218 618008 360704 628385
rect 361089 628508 361139 628732
rect 361523 628508 361575 628732
rect 361089 619534 361575 628508
rect 362010 628699 362496 628770
rect 362010 628475 362055 628699
rect 362439 628475 362496 628699
rect 362010 620980 362496 628475
rect 362010 620494 383337 620980
rect 382851 619658 383337 620494
rect 361089 619048 379241 619534
rect 360218 617522 374744 618008
rect 378755 617971 379241 619048
rect 374258 616445 374744 617522
rect 358816 615836 369845 616322
rect 356365 614551 365990 615037
rect 369359 614999 369845 615836
rect 352226 613265 360609 613751
rect 360123 612028 360609 613265
rect 365504 613072 365990 614551
rect 209899 607175 210159 611719
rect 212223 607175 212399 611719
rect 209899 606979 212399 607175
rect 152609 510212 152634 510668
rect 153810 510212 153837 510668
rect 152609 510169 153837 510212
rect 144145 467018 144193 467314
rect 145449 467018 145521 467314
rect 144145 466948 145521 467018
rect -800 465944 480 466056
rect -800 464872 1188 464874
rect -800 464762 1508 464872
rect 253 464760 1508 464762
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 359161 315293 361661 612028
rect 363819 361386 366319 613072
rect 368397 407710 370897 614999
rect 373136 452031 375636 616445
rect 377553 496436 380053 617971
rect 381890 581162 384390 619658
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 570571 584856 580767 585210
rect 570571 584744 584800 584856
rect 570571 582710 580767 584744
rect 583520 583562 584800 583674
rect 570571 581162 573071 582710
rect 381890 578662 573071 581162
rect 582340 555254 584800 555362
rect 582340 554118 582458 555254
rect 582330 554054 582458 554118
rect 584682 554118 584800 555254
rect 584682 554054 584810 554118
rect 582330 551670 582378 554054
rect 584762 551670 584810 554054
rect 582330 551658 582458 551670
rect 582340 550630 582458 551658
rect 584682 551658 584810 551670
rect 584682 550630 584800 551658
rect 582340 550562 584800 550630
rect 582340 545150 584800 545362
rect 582340 540686 582503 545150
rect 584647 540686 584800 545150
rect 582340 540562 584800 540686
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 377553 495434 581308 496436
rect 377553 495322 584800 495434
rect 377553 493936 581308 495322
rect 583520 494140 584800 494252
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 373136 451012 581762 452031
rect 373136 450900 584800 451012
rect 373136 449531 581762 450900
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 368397 406590 581354 407710
rect 583520 407660 584800 407772
rect 368397 406478 584800 406590
rect 368397 405210 581354 406478
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 363819 360168 580825 361386
rect 583520 361238 584800 361350
rect 363819 360056 584800 360168
rect 363819 358886 580825 360056
rect 583520 358874 584800 358986
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 359161 314946 581320 315293
rect 359161 314834 584800 314946
rect 359161 312793 581320 314834
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 578927 240561 584011 240589
rect 578927 224977 578957 240561
rect 583981 240030 584011 240561
rect 583981 235230 584800 240030
rect 583981 230030 584011 235230
rect 583981 225230 584800 230030
rect 583981 224977 584011 225230
rect 578927 224950 584011 224977
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 151577 584800 151630
rect 578897 151565 584800 151577
rect 578897 136621 578908 151565
rect 583772 146830 584800 151565
rect 583772 141630 583784 146830
rect 583772 136830 584800 141630
rect 583772 136621 583784 136830
rect 578897 136610 583784 136621
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 17558 690841 19942 693225
rect 66218 690836 68522 693220
rect 21901 681731 22845 683875
rect 23057 660647 64001 661237
rect 23057 660133 23065 660647
rect 23065 660133 64001 660647
rect 93859 693936 95763 695840
rect 93870 681813 95694 683877
rect 125008 690380 125952 692284
rect 83766 660820 124070 661465
rect 83766 660204 83777 660820
rect 83777 660204 124070 660820
rect 83766 660201 124070 660204
rect 14463 621651 64607 624595
rect 2674 607097 4978 611721
rect 83169 622046 133393 624590
rect 211682 694007 214066 695751
rect 218739 694913 221043 697297
rect 223943 694942 226247 697326
rect 207618 690349 209922 692333
rect 190393 664818 192857 667282
rect 157083 660495 197707 660499
rect 157083 659479 157087 660495
rect 157087 659479 197703 660495
rect 197703 659479 197707 660495
rect 157083 659475 197707 659479
rect 242750 699652 245214 702116
rect 228987 694956 231291 697340
rect 227301 688638 230725 688661
rect 227301 688117 227305 688638
rect 227305 688117 230721 688638
rect 230721 688117 230725 688638
rect 202809 685269 247113 685278
rect 202809 684733 202813 685269
rect 202813 684734 247109 685269
rect 247109 684734 247113 685269
rect 202813 684733 247033 684734
rect 202809 684094 247033 684733
rect 137770 607191 139754 611815
rect 156516 620746 206820 624090
rect 510307 701813 525571 704677
rect 510467 697733 525571 701813
rect 567893 696734 570357 698718
rect 414582 693939 417046 696403
rect 466738 693939 469202 696403
rect 313064 669246 315528 671710
rect 309412 665676 311876 668140
rect 305196 662188 307660 664652
rect 301243 659173 303707 661637
rect 296908 655858 299372 658322
rect 576304 679186 578288 681650
rect 373478 669246 374822 671710
rect 371791 665676 373135 668140
rect 369976 662188 371320 664652
rect 368202 659173 369546 661637
rect 366163 655858 367507 658322
rect 325573 648381 328037 650845
rect 347669 636730 348053 637114
rect 352237 630050 352701 630274
rect 356376 630031 356840 630255
rect 358827 630053 359291 630277
rect 360271 628385 360655 628609
rect 361139 628508 361523 628732
rect 362055 628475 362439 628699
rect 210159 607175 212223 611719
rect 582458 554054 584682 555254
rect 582378 551670 584762 554054
rect 582458 550630 584682 551670
rect 582503 540686 584647 545150
rect 578957 224977 583981 240561
rect 578908 136621 583772 151565
<< metal4 >>
rect 510305 704683 525574 704717
rect 510305 704677 510461 704683
rect 525417 704677 525574 704683
rect 242731 702122 245233 702135
rect 242731 699646 242744 702122
rect 245220 699646 245233 702122
rect 510305 701813 510307 704677
rect 510305 701789 510467 701813
rect 242731 699633 245233 699646
rect 510465 697733 510467 701789
rect 525571 697733 525574 704677
rect 510465 697727 510781 697733
rect 525417 697727 525574 697733
rect 510465 697693 525574 697727
rect 567874 698718 570376 698737
rect 218687 697340 231368 697368
rect 218687 697326 228987 697340
rect 218687 697297 223943 697326
rect 93805 695840 214125 695904
rect 93805 693936 93859 695840
rect 95763 695751 214125 695840
rect 95763 694007 211682 695751
rect 214066 694007 214125 695751
rect 218687 694913 218739 697297
rect 221043 694942 223943 697297
rect 226247 694956 228987 697326
rect 231291 694956 231368 697340
rect 567874 696734 567893 698718
rect 570357 696734 570376 698718
rect 567874 696716 570376 696734
rect 226247 694942 231368 694956
rect 221043 694913 231368 694942
rect 218687 694868 231368 694913
rect 414563 696409 417065 696422
rect 95763 693936 214125 694007
rect 93805 693889 214125 693936
rect 414563 693933 414576 696409
rect 417052 693933 417065 696409
rect 414563 693920 417065 693933
rect 466719 696409 469221 696422
rect 466719 693933 466732 696409
rect 469208 693933 469221 696409
rect 466719 693920 469221 693933
rect 17498 693225 68630 693269
rect 17498 690841 17558 693225
rect 19942 693220 68630 693225
rect 19942 690841 66218 693220
rect 17498 690836 66218 690841
rect 68522 690836 68630 693220
rect 207590 692349 209951 692356
rect 17498 690769 68630 690836
rect 124977 692333 209951 692349
rect 124977 692284 207618 692333
rect 124977 690380 125008 692284
rect 125952 690380 207618 692284
rect 124977 690349 207618 690380
rect 209922 690349 209951 692333
rect 124977 690334 209951 690349
rect 207590 690327 209951 690334
rect 567875 690311 570375 696716
rect 227276 688661 230751 688665
rect 227276 688507 227301 688661
rect 230725 688507 230751 688661
rect 227276 688271 227295 688507
rect 230731 688271 230751 688507
rect 227276 688117 227301 688271
rect 230725 688117 230751 688271
rect 227276 688114 230751 688117
rect 536686 687811 570375 690311
rect 202779 685278 247143 685292
rect 202779 685235 202809 685278
rect 202733 684094 202809 685235
rect 247113 684734 247143 685278
rect 247033 684710 247143 684734
rect 247033 684094 247110 684710
rect 21910 683907 95867 683939
rect 21891 683877 95867 683907
rect 21891 683875 93870 683877
rect 21891 681731 21901 683875
rect 22845 681813 93870 683875
rect 95694 681813 95867 683877
rect 202733 683308 202883 684094
rect 246959 684081 247110 684094
rect 246959 683308 247109 684081
rect 202733 683217 247109 683308
rect 22845 681731 95867 681813
rect 21891 681710 95867 681731
rect 21891 681700 22855 681710
rect 260437 678032 274962 678175
rect 260437 677902 260541 678032
rect 31160 677834 260541 677902
rect 31160 677668 72152 677834
rect 31049 677609 72152 677668
rect 31049 673213 31133 677609
rect 46409 673213 72152 677609
rect 31049 673154 72152 673213
rect 31160 673118 72152 673154
rect 75268 677819 260541 677834
rect 75268 677707 142945 677819
rect 75268 673311 101969 677707
rect 117565 673311 142945 677707
rect 75268 673118 142945 673311
rect 31160 673103 142945 673118
rect 145421 677775 260541 677819
rect 145421 677662 216598 677775
rect 145421 673266 171414 677662
rect 184770 673266 216598 677662
rect 145421 673103 216598 673266
rect 31160 673059 216598 673103
rect 232194 673059 260541 677775
rect 31160 673035 260541 673059
rect 216578 672994 232215 673035
rect 260437 672036 260541 673035
rect 274857 677902 274962 678032
rect 274857 677825 467817 677902
rect 274857 673109 452357 677825
rect 466993 673109 467817 677825
rect 274857 673035 467817 673109
rect 274857 672036 274962 673035
rect 260437 671893 274962 672036
rect 313045 671728 315547 671729
rect 373474 671728 374826 671729
rect 313045 671710 374835 671728
rect 313045 669246 313064 671710
rect 315528 669246 373478 671710
rect 374822 669246 374835 671710
rect 313045 669228 374835 669246
rect 313045 669227 315547 669228
rect 373474 669227 374826 669228
rect 309393 668158 311895 668159
rect 371787 668158 373139 668159
rect 309393 668140 373148 668158
rect 190376 667299 192875 667306
rect 190376 667282 235517 667299
rect 190376 664818 190393 667282
rect 192857 664818 235517 667282
rect 309393 665676 309412 668140
rect 311876 665676 371791 668140
rect 373135 665676 373148 668140
rect 309393 665658 373148 665676
rect 309393 665657 311895 665658
rect 371787 665657 373139 665658
rect 190376 664799 235517 664818
rect 190376 664795 192875 664799
rect 83765 662744 124085 662834
rect 23042 661749 64017 661882
rect 23042 661270 23091 661749
rect 23041 661237 23091 661270
rect 63967 661270 64017 661749
rect 83765 661488 83807 662744
rect 83764 661465 83807 661488
rect 124043 661465 124085 662744
rect 63967 661237 64018 661270
rect 23041 660133 23057 661237
rect 64001 660133 64018 661237
rect 83764 660201 83766 661465
rect 124070 660201 124085 661465
rect 157083 661364 197702 661420
rect 157083 660503 157114 661364
rect 83764 660179 124085 660201
rect 157082 660499 157114 660503
rect 197670 660503 197702 661364
rect 197670 660499 197709 660503
rect 83764 660178 124072 660179
rect 23041 660100 64018 660133
rect 157082 659475 157083 660499
rect 197707 659475 197709 660499
rect 157082 659471 197709 659475
rect 233017 635570 235517 664799
rect 305177 664670 307679 664671
rect 369972 664670 371324 664671
rect 305177 664652 371333 664670
rect 305177 662188 305196 664652
rect 307660 662188 369976 664652
rect 371320 662188 371333 664652
rect 305177 662170 371333 662188
rect 305177 662169 307679 662170
rect 369972 662169 371324 662170
rect 301224 661655 303726 661656
rect 368198 661655 369550 661656
rect 301224 661637 369559 661655
rect 301224 659173 301243 661637
rect 303707 659173 368202 661637
rect 369546 659173 369559 661637
rect 301224 659155 369559 659173
rect 301224 659154 303726 659155
rect 368198 659154 369550 659155
rect 296889 658340 299391 658341
rect 366159 658340 367511 658341
rect 296889 658322 367520 658340
rect 296889 655858 296908 658322
rect 299372 655858 366163 658322
rect 367507 655858 367520 658322
rect 296889 655840 367520 655858
rect 296889 655839 299391 655840
rect 366159 655839 367511 655840
rect 325554 650863 328056 650864
rect 251036 650845 328065 650863
rect 251036 648381 325573 650845
rect 328037 648381 328065 650845
rect 251036 648363 328065 648381
rect 251036 643769 253536 648363
rect 325554 648362 328056 648363
rect 356670 643894 356990 643930
rect 251036 641269 338266 643769
rect 356670 643658 356712 643894
rect 356948 643763 356990 643894
rect 359056 643894 359376 643930
rect 359056 643763 359098 643894
rect 356948 643658 357847 643763
rect 356670 643636 357847 643658
rect 356670 643622 356990 643636
rect 357720 642897 357847 643636
rect 358200 643658 359098 643763
rect 359334 643658 359376 643894
rect 358200 643636 359376 643658
rect 358200 642897 358327 643636
rect 359056 643622 359376 643636
rect 335766 640142 338266 641269
rect 335766 639692 348716 640142
rect 536686 639819 539186 687811
rect 576286 681668 578307 681669
rect 360315 637525 360607 637553
rect 360315 637289 360343 637525
rect 360579 637289 360607 637525
rect 360315 637262 360607 637289
rect 361033 637515 361327 637566
rect 361033 637279 361062 637515
rect 361298 637279 361327 637515
rect 361033 637228 361327 637279
rect 362102 637532 362396 637583
rect 362102 637296 362131 637532
rect 362367 637296 362396 637532
rect 362102 637245 362396 637296
rect 383342 637319 539186 639819
rect 544840 681650 578307 681668
rect 544840 679186 576304 681650
rect 578288 679186 578307 681650
rect 544840 679168 578307 679186
rect 347635 637147 348087 637148
rect 335766 637114 348087 637147
rect 335766 636730 347669 637114
rect 348053 636730 348087 637114
rect 335766 636697 348087 636730
rect 335766 635570 338266 636697
rect 347635 636696 348087 636697
rect 383342 635788 383892 637319
rect 376970 635579 383892 635788
rect 233017 633070 338266 635570
rect 376994 633304 383892 633513
rect 352335 630282 352605 632949
rect 352235 630274 352703 630282
rect 352235 630050 352237 630274
rect 352701 630050 352703 630274
rect 356477 630263 356747 632977
rect 358930 630285 359200 632879
rect 383342 631773 383892 633304
rect 544840 631773 547340 679168
rect 576286 679167 578307 679168
rect 358825 630277 359293 630285
rect 352235 630043 352703 630050
rect 356374 630255 356842 630263
rect 356374 630031 356376 630255
rect 356840 630031 356842 630255
rect 358825 630053 358827 630277
rect 359291 630053 359293 630277
rect 358825 630046 359293 630053
rect 356374 630024 356842 630031
rect 383342 629273 547340 631773
rect 361131 628738 361531 628772
rect 361131 628732 361213 628738
rect 361449 628732 361531 628738
rect 360263 628615 360663 628649
rect 360263 628609 360345 628615
rect 360581 628609 360663 628615
rect 360263 628385 360271 628609
rect 360655 628385 360663 628609
rect 361131 628508 361139 628732
rect 361523 628508 361531 628732
rect 361131 628502 361213 628508
rect 361449 628502 361531 628508
rect 361131 628468 361531 628502
rect 362047 628705 362447 628739
rect 362047 628699 362129 628705
rect 362365 628699 362447 628705
rect 362047 628475 362055 628699
rect 362439 628475 362447 628699
rect 362047 628469 362129 628475
rect 362365 628469 362447 628475
rect 362047 628435 362447 628469
rect 360263 628379 360345 628385
rect 360581 628379 360663 628385
rect 360263 628345 360663 628379
rect 259670 625130 275302 625270
rect 83049 624683 133410 624733
rect 82973 624631 133488 624683
rect 14426 624595 64645 624620
rect 14426 624437 14463 624595
rect 14337 624377 14463 624437
rect 14337 618061 14391 624377
rect 64607 621651 64645 624595
rect 64227 621626 64645 621651
rect 64227 618061 64282 621626
rect 14337 618001 64282 618061
rect 82973 617995 82992 624631
rect 133468 617995 133488 624631
rect 156499 624090 206837 624129
rect 156499 624087 156516 624090
rect 156376 620746 156516 624087
rect 206820 620746 206837 624090
rect 156376 619257 156528 620746
rect 206684 620708 206837 620746
rect 206684 619257 206836 620708
rect 156376 619144 206836 619257
rect 82973 617893 133488 617995
rect 259670 617214 259688 625130
rect 275284 625028 275302 625130
rect 275284 624590 345528 625028
rect 275284 617634 311401 624590
rect 345237 623908 345528 624590
rect 345237 623829 380589 623908
rect 345237 623593 380249 623829
rect 380485 623593 380589 623829
rect 345237 623509 380589 623593
rect 345237 623273 380249 623509
rect 380485 623273 380589 623509
rect 345237 623189 380589 623273
rect 345237 622953 380249 623189
rect 380485 622953 380589 623189
rect 345237 622869 380589 622953
rect 345237 622633 380249 622869
rect 380485 622633 380589 622869
rect 345237 622549 380589 622633
rect 345237 622313 380249 622549
rect 380485 622313 380589 622549
rect 345237 622229 380589 622313
rect 345237 621993 380249 622229
rect 380485 621993 380589 622229
rect 345237 621915 380589 621993
rect 345237 617634 345528 621915
rect 275284 617272 345528 617634
rect 275284 617214 275302 617272
rect 259670 617074 275302 617214
rect 2575 611815 212044 611907
rect 2575 611721 137770 611815
rect 2575 607097 2674 611721
rect 4978 607191 137770 611721
rect 139754 611734 212044 611815
rect 139754 611719 212246 611734
rect 139754 607191 210159 611719
rect 4978 607175 210159 607191
rect 212223 607175 212246 611719
rect 4978 607160 212246 607175
rect 4978 607097 212044 607160
rect 2575 607040 212044 607097
rect 30038 599270 561785 599316
rect 30038 583994 30289 599270
rect 45885 599167 561785 599270
rect 45885 599156 381236 599167
rect 45885 599110 124972 599156
rect 45885 598950 77177 599110
rect 30038 583674 41489 583994
rect 67325 583674 77177 598950
rect 30038 583514 77177 583674
rect 79653 598838 124972 599110
rect 79653 583514 100792 598838
rect 30038 583445 100792 583514
rect 100668 583242 100792 583445
rect 116388 583560 124972 598838
rect 154648 599109 381236 599156
rect 154648 599011 289763 599109
rect 154648 598789 195952 599011
rect 154648 583833 172492 598789
rect 187768 583833 195952 598789
rect 154648 583735 195952 583833
rect 227868 583735 289763 599011
rect 154648 583560 289763 583735
rect 116388 583513 289763 583560
rect 319439 598624 381236 599109
rect 319439 583988 338634 598624
rect 353910 583988 381236 598624
rect 319439 583571 381236 583988
rect 410912 599148 561785 599167
rect 410912 583571 487943 599148
rect 319439 583552 487943 583571
rect 525619 598751 561785 599148
rect 525619 584115 546218 598751
rect 561174 584115 561785 598751
rect 525619 583552 561785 584115
rect 319439 583513 561785 583552
rect 116388 583445 561785 583513
rect 116388 583242 116512 583445
rect 100668 583221 116512 583242
rect 20619 555772 584769 555900
rect 17921 555625 584769 555772
rect 17921 540349 17943 555625
rect 32899 555515 584769 555625
rect 32899 555414 259906 555515
rect 32899 555334 199833 555414
rect 32899 540378 41075 555334
rect 70751 555197 199833 555334
rect 70751 540561 129115 555197
rect 159111 540561 199833 555197
rect 70751 540458 199833 540561
rect 229829 540559 259906 555414
rect 275182 555513 584769 555515
rect 275182 555434 452190 555513
rect 275182 555159 385288 555434
rect 275182 540559 293931 555159
rect 229829 540523 293931 540559
rect 323927 540798 385288 555159
rect 415284 540798 452190 555434
rect 323927 540523 452190 540798
rect 229829 540458 452190 540523
rect 70751 540378 452190 540458
rect 32899 540349 452190 540378
rect 17921 540237 452190 540349
rect 467466 555254 584769 555513
rect 467466 555225 582458 555254
rect 467466 540589 491316 555225
rect 521952 554054 582458 555225
rect 584682 554119 584769 555254
rect 584682 554054 584801 554119
rect 521952 551670 582378 554054
rect 584762 551670 584801 554054
rect 521952 550630 582458 551670
rect 584682 551657 584801 551670
rect 584682 550630 584769 551657
rect 521952 549950 584769 550630
rect 521952 546246 582340 549950
rect 521952 545150 585071 546246
rect 521952 540686 582503 545150
rect 584647 540686 585071 545150
rect 521952 540589 585071 540686
rect 467466 540237 585071 540589
rect 17921 540202 585071 540237
rect 20619 540029 585071 540202
rect 102586 432558 557291 432965
rect 101051 432468 557291 432558
rect 101051 417512 101088 432468
rect 116364 417832 338922 432468
rect 354198 432093 557291 432468
rect 354198 432002 561038 432093
rect 354198 417832 545733 432002
rect 116364 417512 545733 417832
rect 101051 417422 545733 417512
rect 102586 417366 545733 417422
rect 561009 417366 561038 432002
rect 102586 417276 561038 417366
rect 102586 417094 557291 417276
rect 21612 378918 466454 379014
rect 21612 378829 467213 378918
rect 21612 378665 452175 378829
rect 21612 378616 260096 378665
rect 17721 378460 260096 378616
rect 17721 363504 17733 378460
rect 33009 363504 260096 378460
rect 17721 363389 260096 363504
rect 275052 363553 452175 378665
rect 467131 363553 467213 378829
rect 275052 363464 467213 363553
rect 275052 363389 466454 363464
rect 17721 363349 466454 363389
rect 21612 363143 466454 363349
rect 22911 240605 583937 240685
rect 17911 240590 583937 240605
rect 17911 240561 584002 240590
rect 17911 240491 578957 240561
rect 17911 225215 17985 240491
rect 32621 240343 578957 240491
rect 32621 240321 452145 240343
rect 32621 225365 259905 240321
rect 274861 225387 452145 240321
rect 467421 225387 578957 240343
rect 274861 225365 578957 225387
rect 32621 225215 578957 225365
rect 17911 225102 578957 225215
rect 22911 225078 578957 225102
rect 563330 224977 578957 225078
rect 583981 224977 584002 240561
rect 563330 224949 584002 224977
rect 563330 224854 583937 224949
rect 100326 151638 584154 151892
rect 100326 151590 545507 151638
rect 100326 136634 100611 151590
rect 116527 151535 545507 151590
rect 116527 136634 338714 151535
rect 100326 136579 338714 136634
rect 354310 136682 545507 151535
rect 561423 151565 584154 151638
rect 561423 136682 578908 151565
rect 354310 136621 578908 136682
rect 583772 136621 584154 151565
rect 354310 136579 584154 136621
rect 100326 136443 584154 136579
<< via4 >>
rect 510461 704677 525417 704683
rect 242744 702116 245220 702122
rect 242744 699652 242750 702116
rect 242750 699652 245214 702116
rect 245214 699652 245220 702116
rect 242744 699646 245220 699652
rect 510461 701887 525417 704677
rect 510781 697733 525417 701887
rect 510781 697727 525417 697733
rect 414576 696403 417052 696409
rect 414576 693939 414582 696403
rect 414582 693939 417046 696403
rect 417046 693939 417052 696403
rect 414576 693933 417052 693939
rect 466732 696403 469208 696409
rect 466732 693939 466738 696403
rect 466738 693939 469202 696403
rect 469202 693939 469208 696403
rect 466732 693933 469208 693939
rect 227295 688271 227301 688507
rect 227301 688271 227531 688507
rect 227615 688271 227851 688507
rect 227935 688271 228171 688507
rect 228255 688271 228491 688507
rect 228575 688271 228811 688507
rect 228895 688271 229131 688507
rect 229215 688271 229451 688507
rect 229535 688271 229771 688507
rect 229855 688271 230091 688507
rect 230175 688271 230411 688507
rect 230495 688271 230725 688507
rect 230725 688271 230731 688507
rect 202883 684094 246959 685144
rect 202883 683308 246959 684094
rect 31133 673213 46409 677609
rect 72152 673118 75268 677834
rect 101969 673311 117565 677707
rect 142945 673103 145421 677819
rect 171414 673266 184770 677662
rect 216598 673059 232194 677775
rect 260541 672036 274857 678032
rect 452357 673109 466993 677825
rect 23091 661237 63967 661749
rect 83807 661465 124043 662744
rect 23091 660233 63967 661237
rect 83807 660268 124043 661465
rect 157114 660499 197670 661364
rect 157114 659528 197670 660499
rect 356712 643658 356948 643894
rect 359098 643658 359334 643894
rect 360343 637289 360579 637525
rect 361062 637279 361298 637515
rect 362131 637296 362367 637532
rect 361213 628732 361449 628738
rect 360345 628609 360581 628615
rect 360345 628385 360581 628609
rect 361213 628508 361449 628732
rect 361213 628502 361449 628508
rect 362129 628699 362365 628705
rect 362129 628475 362365 628699
rect 362129 628469 362365 628475
rect 360345 628379 360581 628385
rect 14391 621651 14463 624377
rect 14463 621651 64227 624377
rect 14391 618061 64227 621651
rect 82992 624590 133468 624631
rect 82992 622046 83169 624590
rect 83169 622046 133393 624590
rect 133393 622046 133468 624590
rect 82992 617995 133468 622046
rect 156528 620746 206684 623973
rect 156528 619257 206684 620746
rect 259688 617214 275284 625130
rect 311401 617634 345237 624590
rect 380249 623593 380485 623829
rect 380249 623273 380485 623509
rect 380249 622953 380485 623189
rect 380249 622633 380485 622869
rect 380249 622313 380485 622549
rect 380249 621993 380485 622229
rect 30289 598950 45885 599270
rect 30289 583994 67325 598950
rect 41489 583674 67325 583994
rect 77177 583514 79653 599110
rect 100792 583242 116388 598838
rect 124972 583560 154648 599156
rect 172492 583833 187768 598789
rect 195952 583735 227868 599011
rect 289763 583513 319439 599109
rect 338634 583988 353910 598624
rect 381236 583571 410912 599167
rect 487943 583552 525619 599148
rect 546218 584115 561174 598751
rect 17943 540349 32899 555625
rect 41075 540378 70751 555334
rect 129115 540561 159111 555197
rect 199833 540458 229829 555414
rect 259906 540559 275182 555515
rect 293931 540523 323927 555159
rect 385288 540798 415284 555434
rect 452190 540237 467466 555513
rect 491316 540589 521952 555225
rect 101088 417512 116364 432468
rect 338922 417832 354198 432468
rect 545733 417366 561009 432002
rect 17733 363504 33009 378460
rect 260096 363389 275052 378665
rect 452175 363553 467131 378829
rect 17985 225215 32621 240491
rect 259905 225365 274861 240321
rect 452145 225387 467421 240343
rect 100611 136634 116527 151590
rect 338714 136579 354310 151535
rect 545507 136682 561423 151638
<< metal5 >>
rect 510282 704683 525597 704740
rect 510282 703705 510461 704683
rect 242708 702122 245256 702158
rect 242708 699646 242744 702122
rect 245220 699646 245256 702122
rect 242708 699610 245256 699646
rect 510173 701887 510461 703705
rect 525417 703705 525597 704683
rect 242732 693377 245232 699610
rect 510173 697727 510781 701887
rect 525417 697727 525839 703705
rect 414540 696421 417088 696445
rect 466696 696421 469244 696445
rect 414540 696409 436162 696421
rect 414540 693933 414576 696409
rect 417052 693933 436162 696409
rect 414540 693921 436162 693933
rect 414540 693897 417088 693921
rect 227790 690877 245232 693377
rect 227790 688688 230290 690877
rect 433662 690218 436162 693921
rect 227253 688507 230774 688688
rect 227253 688271 227295 688507
rect 227531 688271 227615 688507
rect 227851 688271 227935 688507
rect 228171 688271 228255 688507
rect 228491 688271 228575 688507
rect 228811 688271 228895 688507
rect 229131 688271 229215 688507
rect 229451 688271 229535 688507
rect 229771 688271 229855 688507
rect 230091 688271 230175 688507
rect 230411 688271 230495 688507
rect 230731 688271 230774 688507
rect 227253 688091 230774 688271
rect 352750 687718 436162 690218
rect 441224 696409 469244 696421
rect 441224 693933 466732 696409
rect 469208 693933 469244 696409
rect 441224 693921 469244 693933
rect 202709 685144 247133 685259
rect 202709 683308 202883 685144
rect 246959 683308 247133 685144
rect 202709 683193 247133 683308
rect 30960 677609 46833 678350
rect 30960 673213 31133 677609
rect 46409 673213 46833 677609
rect 30960 661906 46833 673213
rect 72119 677834 75301 677881
rect 72119 673118 72152 677834
rect 75268 677536 75301 677834
rect 142912 677819 145454 677900
rect 216581 677865 232247 683193
rect 101944 677707 117591 677810
rect 75268 673118 75313 677536
rect 101944 677524 101969 677707
rect 72119 673072 75313 673118
rect 23018 661749 64041 661906
rect 23018 660233 23091 661749
rect 63967 660233 64041 661749
rect 23018 660077 64041 660233
rect 14313 624377 64306 624461
rect 14313 618061 14391 624377
rect 64227 618061 64306 624377
rect 14313 617977 64306 618061
rect 30017 599270 46173 617977
rect 72165 615148 75313 673072
rect 101864 673311 101969 677524
rect 117565 677524 117591 677707
rect 142912 677705 142945 677819
rect 117565 673311 117672 677524
rect 77216 613098 79845 671573
rect 101864 662858 117672 673311
rect 142885 673103 142945 677705
rect 145421 677705 145454 677819
rect 145421 673103 145500 677705
rect 171296 677662 184889 677842
rect 171296 677636 171414 677662
rect 83741 662744 124109 662858
rect 83741 660268 83807 662744
rect 124043 660268 124109 662744
rect 83741 660155 124109 660268
rect 83025 624707 133434 624757
rect 82949 624631 133512 624707
rect 82949 617995 82992 624631
rect 133468 617995 133512 624631
rect 82949 617869 133512 617995
rect 30017 586019 30289 599270
rect 45885 599169 46173 599270
rect 51497 599196 53807 599338
rect 58426 599196 60736 599292
rect 65356 599196 67666 599323
rect 51497 599169 67666 599196
rect 45885 598950 67666 599169
rect 30156 583994 30289 586019
rect 30156 583677 41489 583994
rect 36223 560658 38615 583677
rect 41423 583674 41489 583677
rect 67325 583674 67666 598950
rect 41423 583639 67666 583674
rect 44501 581203 46811 583639
rect 51497 581259 53807 583639
rect 45425 580076 45745 581203
rect 52369 580076 52689 581259
rect 58426 581098 60736 583639
rect 65356 581205 67666 583639
rect 77058 599110 79845 613098
rect 77058 583524 77177 599110
rect 77059 583514 77177 583524
rect 79653 583612 79845 599110
rect 100463 598838 116619 617869
rect 142885 615246 145500 673103
rect 171295 673266 171414 677636
rect 184770 673266 184889 677662
rect 171295 673086 184889 673266
rect 216554 677775 232247 677865
rect 79653 583514 79771 583612
rect 77059 583474 79771 583514
rect 100463 583242 100792 598838
rect 116388 583242 116619 598838
rect 59313 580076 59633 581098
rect 66257 580076 66577 581205
rect 17569 555625 33235 556317
rect 17569 540349 17943 555625
rect 32899 540349 33235 555625
rect 17569 378460 33235 540349
rect 40864 555438 43451 578397
rect 48022 555438 50609 578656
rect 54834 555438 57421 578570
rect 61819 555438 64406 578052
rect 68545 555438 71132 578483
rect 40864 555334 71132 555438
rect 40864 540378 41075 555334
rect 70751 540378 71132 555334
rect 40864 540274 71132 540378
rect 40864 540137 43451 540274
rect 48022 540113 50609 540274
rect 54834 540113 57421 540274
rect 61819 540137 64406 540274
rect 68545 540212 71132 540274
rect 17569 363504 17733 378460
rect 33009 363504 33235 378460
rect 17569 240491 33235 363504
rect 17569 225215 17985 240491
rect 32621 225215 33235 240491
rect 17569 224794 33235 225215
rect 100463 432468 116619 583242
rect 124759 599200 126962 599322
rect 147647 599200 151189 672301
rect 171295 661444 184887 673086
rect 216554 673059 216598 677775
rect 232194 673059 232247 677775
rect 216554 673051 232247 673059
rect 259666 678032 275332 678276
rect 216554 672970 232239 673051
rect 157059 661364 197726 661444
rect 157059 659528 157114 661364
rect 197670 659528 197726 661364
rect 157059 659448 197726 659528
rect 156352 624096 206860 624111
rect 156352 623973 207124 624096
rect 156352 619257 156528 623973
rect 206684 619257 207124 623973
rect 156352 619120 207124 619257
rect 154493 599200 154813 599217
rect 124759 599156 154813 599200
rect 124759 583560 124972 599156
rect 154648 583560 154813 599156
rect 172171 598789 188327 619120
rect 218723 615607 222084 672970
rect 259666 672036 260541 678032
rect 274857 672036 275332 678032
rect 223844 599042 227386 658283
rect 259666 625294 275332 672036
rect 352750 647598 355250 687718
rect 441224 684427 443724 693921
rect 466696 693897 469244 693921
rect 360796 681927 443724 684427
rect 360796 647598 363296 681927
rect 352750 647048 356990 647598
rect 356670 643954 356990 647048
rect 359056 647048 363296 647598
rect 451976 677825 467642 678029
rect 451976 673109 452357 677825
rect 466993 673109 467642 677825
rect 359056 643954 359376 647048
rect 356646 643894 357014 643954
rect 356646 643658 356712 643894
rect 356948 643658 357014 643894
rect 356646 643598 357014 643658
rect 359032 643894 359400 643954
rect 359032 643658 359098 643894
rect 359334 643658 359400 643894
rect 359032 643598 359400 643658
rect 360291 637525 360631 637577
rect 360291 637289 360343 637525
rect 360579 637427 360631 637525
rect 361009 637515 361351 637590
rect 360579 637289 360633 637427
rect 259646 625130 275332 625294
rect 259646 617214 259688 625130
rect 275284 617214 275332 625130
rect 344840 624668 345283 631382
rect 346785 627046 347228 631405
rect 360291 628672 360633 637289
rect 361009 637279 361062 637515
rect 361298 637279 361351 637515
rect 361009 636893 361351 637279
rect 362078 637532 362420 637607
rect 362078 637296 362131 637532
rect 362367 637296 362420 637532
rect 361009 628795 361344 636893
rect 361009 628738 361554 628795
rect 362078 628762 362420 637296
rect 360240 628615 360686 628672
rect 360240 628379 360345 628615
rect 360581 628379 360686 628615
rect 361009 628502 361213 628738
rect 361449 628502 361554 628738
rect 361009 628473 361554 628502
rect 361108 628445 361554 628473
rect 362024 628705 362470 628762
rect 362024 628469 362129 628705
rect 362365 628469 362470 628705
rect 362024 628412 362470 628469
rect 360240 628322 360686 628379
rect 378201 627046 378644 630294
rect 346785 625053 378644 627046
rect 311256 624590 345382 624668
rect 311256 617634 311401 624590
rect 345237 617634 345382 624590
rect 311256 617556 345382 617634
rect 259646 617050 275332 617214
rect 195827 599011 227994 599042
rect 195827 598960 195952 599011
rect 172171 583913 172492 598789
rect 172445 583833 172492 583913
rect 187768 583913 188327 598789
rect 187768 583833 187815 583913
rect 172445 583650 187815 583833
rect 195244 583735 195952 598960
rect 227868 583735 227994 599011
rect 195244 583705 227994 583735
rect 124759 583523 154813 583560
rect 124759 560338 126962 583523
rect 133661 579201 133981 583523
rect 140605 579201 140925 583523
rect 147549 583483 151122 583523
rect 147549 578864 147869 583483
rect 154493 579201 154813 583523
rect 195244 579563 197447 583705
rect 195244 579361 197522 579563
rect 128823 555375 131710 577101
rect 135608 555375 138495 576885
rect 143114 555375 146001 576957
rect 149754 555375 152641 577029
rect 156683 555375 159570 576740
rect 195244 573243 197447 579361
rect 197480 573243 197522 579361
rect 204146 579361 204466 583705
rect 197842 579262 203810 579286
rect 197842 573342 197866 579262
rect 199308 573342 202195 577261
rect 203786 573342 203810 579262
rect 197842 573318 203810 573342
rect 195244 572839 197522 573243
rect 195244 566721 197447 572839
rect 197480 566721 197522 572839
rect 199308 572764 202195 573318
rect 204146 573243 204188 579361
rect 204424 573243 204466 579361
rect 211090 579361 211410 583705
rect 204786 579262 210754 579286
rect 204786 573342 204810 579262
rect 206093 573342 208980 577045
rect 210730 573342 210754 579262
rect 204786 573318 210754 573342
rect 204146 572839 204466 573243
rect 197842 572740 203810 572764
rect 197842 566820 197866 572740
rect 199308 566820 202195 572740
rect 203786 566820 203810 572740
rect 197842 566796 203810 566820
rect 195244 566317 197522 566721
rect 195244 560199 197447 566317
rect 197480 560199 197522 566317
rect 199308 566242 202195 566796
rect 204146 566721 204188 572839
rect 204424 566721 204466 572839
rect 206093 572764 208980 573318
rect 211090 573243 211132 579361
rect 211368 573243 211410 579361
rect 211730 579262 216581 579286
rect 211730 573342 211754 579262
rect 218034 579243 218354 583705
rect 224978 579243 225298 583705
rect 213599 573342 216486 577117
rect 211730 573318 216581 573342
rect 211090 572839 211410 573243
rect 204786 572740 210754 572764
rect 204786 566820 204810 572740
rect 206093 566820 208980 572740
rect 210730 566820 210754 572740
rect 204786 566796 210754 566820
rect 204146 566317 204466 566721
rect 197842 566218 203810 566242
rect 197842 560298 197866 566218
rect 199308 560298 202195 566218
rect 203786 560298 203810 566218
rect 197842 560274 203810 560298
rect 195244 560051 197522 560199
rect 197202 559997 197522 560051
rect 128823 555197 159570 555375
rect 128823 540561 129115 555197
rect 159111 540561 159570 555197
rect 128823 540383 159570 540561
rect 199308 555488 202195 560274
rect 204146 560199 204188 566317
rect 204424 560199 204466 566317
rect 206093 566242 208980 566796
rect 211090 566721 211132 572839
rect 211368 566721 211410 572839
rect 213599 572764 216486 573318
rect 211730 572740 216581 572764
rect 211730 566820 211754 572740
rect 213599 566820 216486 572740
rect 211730 566796 216581 566820
rect 211090 566317 211410 566721
rect 204786 566218 210754 566242
rect 204786 560298 204810 566218
rect 206093 560298 208980 566218
rect 210730 560298 210754 566218
rect 204786 560274 210754 560298
rect 204146 559997 204466 560199
rect 206093 555488 208980 560274
rect 211090 560199 211132 566317
rect 211368 560199 211410 566317
rect 213599 566242 216486 566796
rect 211730 566218 216581 566242
rect 211730 560298 211754 566218
rect 213599 560298 216486 566218
rect 211730 560274 216581 560298
rect 211090 559997 211410 560199
rect 213599 555488 216486 560274
rect 220132 555488 223019 578371
rect 227397 555488 230284 578371
rect 199308 555414 230284 555488
rect 199308 540458 199833 555414
rect 229829 540458 230284 555414
rect 199308 540415 230284 540458
rect 259666 555515 275332 617050
rect 312320 604344 315940 617556
rect 319399 604291 323019 617556
rect 326025 604364 329645 617556
rect 333307 604619 336927 617556
rect 340152 604546 343772 617556
rect 346785 615384 354541 625053
rect 380146 623932 380589 631171
rect 380122 623829 380613 623932
rect 380122 623593 380249 623829
rect 380485 623593 380613 623829
rect 380122 623509 380613 623593
rect 380122 623273 380249 623509
rect 380485 623273 380613 623509
rect 380122 623189 380613 623273
rect 380122 622953 380249 623189
rect 380485 622953 380613 623189
rect 380122 622869 380613 622953
rect 380122 622633 380249 622869
rect 380485 622633 380613 622869
rect 380122 622549 380613 622633
rect 380122 622313 380249 622549
rect 380485 622313 380613 622549
rect 380122 622229 380613 622313
rect 380122 621993 380249 622229
rect 380485 621993 380613 622229
rect 380122 621891 380613 621993
rect 345371 602316 354541 615384
rect 317349 600961 317669 602316
rect 324293 600961 324613 602316
rect 331237 600961 331557 602316
rect 338181 600961 338501 602316
rect 345125 600961 354541 602316
rect 317349 600926 354541 600961
rect 289452 599150 291655 599152
rect 317078 599150 354541 600926
rect 289452 599109 354541 599150
rect 289452 583513 289763 599109
rect 319439 598624 354541 599109
rect 381102 599167 411047 599208
rect 381102 598681 381236 599167
rect 319439 598383 338634 598624
rect 319439 583513 319574 598383
rect 338578 597776 338634 598383
rect 289452 583473 319574 583513
rect 338385 583988 338634 597776
rect 353910 583988 354541 598624
rect 289452 579107 291655 583473
rect 289452 578905 291730 579107
rect 289452 572787 291655 578905
rect 291688 572787 291730 578905
rect 298354 578905 298674 583473
rect 292050 578806 298018 578830
rect 292050 572886 292074 578806
rect 293516 572886 296403 576805
rect 297994 572886 298018 578806
rect 292050 572862 298018 572886
rect 289452 572383 291730 572787
rect 289452 566265 291655 572383
rect 291688 566265 291730 572383
rect 293516 572308 296403 572862
rect 298354 572787 298396 578905
rect 298632 572787 298674 578905
rect 305298 578905 305618 583473
rect 298994 578806 304962 578830
rect 298994 572886 299018 578806
rect 300301 572886 303188 576589
rect 304938 572886 304962 578806
rect 298994 572862 304962 572886
rect 298354 572383 298674 572787
rect 292050 572284 298018 572308
rect 292050 566364 292074 572284
rect 293516 566364 296403 572284
rect 297994 566364 298018 572284
rect 292050 566340 298018 566364
rect 289452 565861 291730 566265
rect 289452 560042 291655 565861
rect 291410 559743 291452 560042
rect 291688 559743 291730 565861
rect 293516 565786 296403 566340
rect 298354 566265 298396 572383
rect 298632 566265 298674 572383
rect 300301 572308 303188 572862
rect 305298 572787 305340 578905
rect 305576 572787 305618 578905
rect 312242 578905 312562 583473
rect 305938 578806 311906 578830
rect 305938 572886 305962 578806
rect 307807 572886 310694 576661
rect 311882 572886 311906 578806
rect 305938 572862 311906 572886
rect 305298 572383 305618 572787
rect 298994 572284 304962 572308
rect 298994 566364 299018 572284
rect 300301 566364 303188 572284
rect 304938 566364 304962 572284
rect 298994 566340 304962 566364
rect 298354 565861 298674 566265
rect 292050 565762 298018 565786
rect 292050 559842 292074 565762
rect 293516 559842 296403 565762
rect 297994 559842 298018 565762
rect 292050 559818 298018 559842
rect 291410 559541 291730 559743
rect 259666 540559 259906 555515
rect 275182 540559 275332 555515
rect 199671 540385 229991 540415
rect 128823 540159 131710 540383
rect 135608 540308 138495 540383
rect 149754 540308 152641 540383
rect 156683 540308 159570 540383
rect 100463 417512 101088 432468
rect 116364 417512 116619 432468
rect 100463 151590 116619 417512
rect 259666 378665 275332 540559
rect 293516 555337 296403 559818
rect 298354 559743 298396 565861
rect 298632 559743 298674 565861
rect 300301 565786 303188 566340
rect 305298 566265 305340 572383
rect 305576 566265 305618 572383
rect 307807 572308 310694 572862
rect 312242 572787 312284 578905
rect 312520 572787 312562 578905
rect 319186 578905 319506 583473
rect 312882 578806 318850 578830
rect 312882 572886 312906 578806
rect 314447 572886 317334 576733
rect 318826 572886 318850 578806
rect 312882 572862 318850 572886
rect 312242 572383 312562 572787
rect 305938 572284 311906 572308
rect 305938 566364 305962 572284
rect 307807 566364 310694 572284
rect 311882 566364 311906 572284
rect 305938 566340 311906 566364
rect 305298 565861 305618 566265
rect 298994 565762 304962 565786
rect 298994 559842 299018 565762
rect 300301 559842 303188 565762
rect 304938 559842 304962 565762
rect 298994 559818 304962 559842
rect 298354 559541 298674 559743
rect 300301 555337 303188 559818
rect 305298 559743 305340 565861
rect 305576 559743 305618 565861
rect 307807 565786 310694 566340
rect 312242 566265 312284 572383
rect 312520 566265 312562 572383
rect 314447 572308 317334 572862
rect 319186 572787 319228 578905
rect 319464 572787 319506 578905
rect 319826 578806 325794 578830
rect 319826 572886 319850 578806
rect 321376 572886 324263 576444
rect 325770 572886 325794 578806
rect 319826 572862 325794 572886
rect 319186 572383 319506 572787
rect 312882 572284 318850 572308
rect 312882 566364 312906 572284
rect 314447 566364 317334 572284
rect 318826 566364 318850 572284
rect 312882 566340 318850 566364
rect 312242 565861 312562 566265
rect 305938 565762 311906 565786
rect 305938 559842 305962 565762
rect 307807 559842 310694 565762
rect 311882 559842 311906 565762
rect 305938 559818 311906 559842
rect 305298 559541 305618 559743
rect 307807 555337 310694 559818
rect 312242 559743 312284 565861
rect 312520 559743 312562 565861
rect 314447 565786 317334 566340
rect 319186 566265 319228 572383
rect 319464 566265 319506 572383
rect 321376 572308 324263 572862
rect 319826 572284 325794 572308
rect 319826 566364 319850 572284
rect 321376 566364 324263 572284
rect 325770 566364 325794 572284
rect 319826 566340 325794 566364
rect 319186 565861 319506 566265
rect 312882 565762 318850 565786
rect 312882 559842 312906 565762
rect 314447 559842 317334 565762
rect 318826 559842 318850 565762
rect 312882 559818 318850 559842
rect 312242 559541 312562 559743
rect 314447 555337 317334 559818
rect 319186 559743 319228 565861
rect 319464 559743 319506 565861
rect 321376 565786 324263 566340
rect 319826 565762 325794 565786
rect 319826 559842 319850 565762
rect 321376 559842 324263 565762
rect 325770 559842 325794 565762
rect 319826 559818 325794 559842
rect 319186 559541 319506 559743
rect 321376 555337 324263 559818
rect 293516 555159 324263 555337
rect 293516 540523 293931 555159
rect 323927 540523 324263 555159
rect 293516 540392 324263 540523
rect 293516 540345 324092 540392
rect 293516 540198 296403 540345
rect 314447 540295 317334 540345
rect 259666 363389 260096 378665
rect 275052 363389 275332 378665
rect 259666 240321 275332 363389
rect 259666 225941 259905 240321
rect 259731 225365 259905 225941
rect 274861 225941 275332 240321
rect 338385 432468 354541 583988
rect 380930 583571 381236 598681
rect 410912 583571 411047 599167
rect 380930 583531 411047 583571
rect 380930 579563 383133 583531
rect 380930 579361 383208 579563
rect 380930 573243 383133 579361
rect 383166 573243 383208 579361
rect 389832 579361 390152 583531
rect 383528 579262 389496 579286
rect 383528 573342 383552 579262
rect 384994 573342 387881 577261
rect 389472 573342 389496 579262
rect 383528 573318 389496 573342
rect 380930 572839 383208 573243
rect 380930 566721 383133 572839
rect 383166 566721 383208 572839
rect 384994 572764 387881 573318
rect 389832 573243 389874 579361
rect 390110 573243 390152 579361
rect 396776 579361 397096 583531
rect 390472 579262 396440 579286
rect 390472 573342 390496 579262
rect 391779 573342 394666 577045
rect 396416 573342 396440 579262
rect 390472 573318 396440 573342
rect 389832 572839 390152 573243
rect 383528 572740 389496 572764
rect 383528 566820 383552 572740
rect 384994 566820 387881 572740
rect 389472 566820 389496 572740
rect 383528 566796 389496 566820
rect 380930 566317 383208 566721
rect 380930 560498 383133 566317
rect 382888 560199 382930 560498
rect 383166 560199 383208 566317
rect 384994 566242 387881 566796
rect 389832 566721 389874 572839
rect 390110 566721 390152 572839
rect 391779 572764 394666 573318
rect 396776 573243 396818 579361
rect 397054 573243 397096 579361
rect 403720 579361 404040 583531
rect 397416 579262 403384 579286
rect 397416 573342 397440 579262
rect 399285 573342 402172 577117
rect 403360 573342 403384 579262
rect 397416 573318 403384 573342
rect 396776 572839 397096 573243
rect 390472 572740 396440 572764
rect 390472 566820 390496 572740
rect 391779 566820 394666 572740
rect 396416 566820 396440 572740
rect 390472 566796 396440 566820
rect 389832 566317 390152 566721
rect 383528 566218 389496 566242
rect 383528 560298 383552 566218
rect 384994 560298 387881 566218
rect 389472 560298 389496 566218
rect 383528 560274 389496 560298
rect 382888 559997 383208 560199
rect 384994 555612 387881 560274
rect 389832 560199 389874 566317
rect 390110 560199 390152 566317
rect 391779 566242 394666 566796
rect 396776 566721 396818 572839
rect 397054 566721 397096 572839
rect 399285 572764 402172 573318
rect 403720 573243 403762 579361
rect 403998 573243 404040 579361
rect 410664 579361 410984 583531
rect 404360 579262 410328 579286
rect 404360 573342 404384 579262
rect 405925 573342 408812 577189
rect 410304 573342 410328 579262
rect 404360 573318 410328 573342
rect 403720 572839 404040 573243
rect 397416 572740 403384 572764
rect 397416 566820 397440 572740
rect 399285 566820 402172 572740
rect 403360 566820 403384 572740
rect 397416 566796 403384 566820
rect 396776 566317 397096 566721
rect 390472 566218 396440 566242
rect 390472 560298 390496 566218
rect 391779 560298 394666 566218
rect 396416 560298 396440 566218
rect 390472 560274 396440 560298
rect 389832 559997 390152 560199
rect 391779 555612 394666 560274
rect 396776 560199 396818 566317
rect 397054 560199 397096 566317
rect 399285 566242 402172 566796
rect 403720 566721 403762 572839
rect 403998 566721 404040 572839
rect 405925 572764 408812 573318
rect 410664 573243 410706 579361
rect 410942 573243 410984 579361
rect 411304 579262 417272 579286
rect 411304 573342 411328 579262
rect 412854 573342 415741 576900
rect 417248 573342 417272 579262
rect 411304 573318 417272 573342
rect 410664 572839 410984 573243
rect 404360 572740 410328 572764
rect 404360 566820 404384 572740
rect 405925 566820 408812 572740
rect 410304 566820 410328 572740
rect 404360 566796 410328 566820
rect 403720 566317 404040 566721
rect 397416 566218 403384 566242
rect 397416 560298 397440 566218
rect 399285 560298 402172 566218
rect 403360 560298 403384 566218
rect 397416 560274 403384 560298
rect 396776 559997 397096 560199
rect 399285 555612 402172 560274
rect 403720 560199 403762 566317
rect 403998 560199 404040 566317
rect 405925 566242 408812 566796
rect 410664 566721 410706 572839
rect 410942 566721 410984 572839
rect 412854 572764 415741 573318
rect 411304 572740 417272 572764
rect 411304 566820 411328 572740
rect 412854 566820 415741 572740
rect 417248 566820 417272 572740
rect 411304 566796 417272 566820
rect 410664 566317 410984 566721
rect 404360 566218 410328 566242
rect 404360 560298 404384 566218
rect 405925 560298 408812 566218
rect 410304 560298 410328 566218
rect 404360 560274 410328 560298
rect 403720 559997 404040 560199
rect 405925 555612 408812 560274
rect 410664 560199 410706 566317
rect 410942 560199 410984 566317
rect 412854 566242 415741 566796
rect 411304 566218 417272 566242
rect 411304 560298 411328 566218
rect 412854 560298 415741 566218
rect 417248 560298 417272 566218
rect 411304 560274 417272 560298
rect 410664 559997 410984 560199
rect 412854 555612 415741 560274
rect 384994 555434 415741 555612
rect 384994 540798 385288 555434
rect 415284 540798 415741 555434
rect 384994 540633 415741 540798
rect 385124 540620 415741 540633
rect 391779 540524 394666 540620
rect 412854 540415 415741 540620
rect 451976 555513 467642 673109
rect 510173 599189 525839 697727
rect 487908 599148 525839 599189
rect 487908 598849 487943 599148
rect 487426 583552 487943 598849
rect 525619 583552 525839 599148
rect 546152 598751 561241 598824
rect 546152 598734 546218 598751
rect 487426 583512 525839 583552
rect 487426 580018 489629 583512
rect 487426 579816 489704 580018
rect 487426 573698 489629 579816
rect 489662 573698 489704 579816
rect 496328 579816 496648 583512
rect 490024 579717 495992 579741
rect 490024 573797 490048 579717
rect 491490 573797 494377 577716
rect 495968 573797 495992 579717
rect 490024 573773 495992 573797
rect 487426 573294 489704 573698
rect 487426 567176 489629 573294
rect 489662 567176 489704 573294
rect 491490 573219 494377 573773
rect 496328 573698 496370 579816
rect 496606 573698 496648 579816
rect 503272 579816 503592 583512
rect 510173 583472 525839 583512
rect 545384 584115 546218 598734
rect 561174 598734 561241 598751
rect 561174 584115 561540 598734
rect 496968 579717 502936 579741
rect 496968 573797 496992 579717
rect 498275 573797 501162 577500
rect 502912 573797 502936 579717
rect 496968 573773 502936 573797
rect 496328 573294 496648 573698
rect 490024 573195 495992 573219
rect 490024 567275 490048 573195
rect 491490 567275 494377 573195
rect 495968 567275 495992 573195
rect 490024 567251 495992 567275
rect 487426 566772 489704 567176
rect 487426 560953 489629 566772
rect 489384 560654 489426 560953
rect 489662 560654 489704 566772
rect 491490 566697 494377 567251
rect 496328 567176 496370 573294
rect 496606 567176 496648 573294
rect 498275 573219 501162 573773
rect 503272 573698 503314 579816
rect 503550 573698 503592 579816
rect 510216 579816 510536 583472
rect 503912 579717 509880 579741
rect 503912 573797 503936 579717
rect 505781 573797 508668 577572
rect 509856 573797 509880 579717
rect 503912 573773 509880 573797
rect 503272 573294 503592 573698
rect 496968 573195 502936 573219
rect 496968 567275 496992 573195
rect 498275 567275 501162 573195
rect 502912 567275 502936 573195
rect 496968 567251 502936 567275
rect 496328 566772 496648 567176
rect 490024 566673 495992 566697
rect 490024 560753 490048 566673
rect 491490 560753 494377 566673
rect 495968 560753 495992 566673
rect 490024 560729 495992 560753
rect 489384 560452 489704 560654
rect 338385 417832 338922 432468
rect 354198 417832 354541 432468
rect 274861 225365 275035 225941
rect 259731 225236 275035 225365
rect 100463 136634 100611 151590
rect 116527 136634 116619 151590
rect 338385 151535 354541 417832
rect 451976 540237 452190 555513
rect 467466 540237 467642 555513
rect 491490 555373 494377 560729
rect 496328 560654 496370 566772
rect 496606 560654 496648 566772
rect 498275 566697 501162 567251
rect 503272 567176 503314 573294
rect 503550 567176 503592 573294
rect 505781 573219 508668 573773
rect 510216 573698 510258 579816
rect 510494 573698 510536 579816
rect 517160 579816 517480 583472
rect 510856 579717 516824 579741
rect 510856 573797 510880 579717
rect 512421 573797 515308 577644
rect 516800 573797 516824 579717
rect 510856 573773 516824 573797
rect 510216 573294 510536 573698
rect 503912 573195 509880 573219
rect 503912 567275 503936 573195
rect 505781 567275 508668 573195
rect 509856 567275 509880 573195
rect 503912 567251 509880 567275
rect 503272 566772 503592 567176
rect 496968 566673 502936 566697
rect 496968 560753 496992 566673
rect 498275 560753 501162 566673
rect 502912 560753 502936 566673
rect 496968 560729 502936 560753
rect 496328 560452 496648 560654
rect 498275 555373 501162 560729
rect 503272 560654 503314 566772
rect 503550 560654 503592 566772
rect 505781 566697 508668 567251
rect 510216 567176 510258 573294
rect 510494 567176 510536 573294
rect 512421 573219 515308 573773
rect 517160 573698 517202 579816
rect 517438 573698 517480 579816
rect 517800 579717 523768 579741
rect 517800 573797 517824 579717
rect 519350 573797 522237 577355
rect 523744 573797 523768 579717
rect 517800 573773 523768 573797
rect 517160 573294 517480 573698
rect 510856 573195 516824 573219
rect 510856 567275 510880 573195
rect 512421 567275 515308 573195
rect 516800 567275 516824 573195
rect 510856 567251 516824 567275
rect 510216 566772 510536 567176
rect 503912 566673 509880 566697
rect 503912 560753 503936 566673
rect 505781 560753 508668 566673
rect 509856 560753 509880 566673
rect 503912 560729 509880 560753
rect 503272 560452 503592 560654
rect 505781 555373 508668 560729
rect 510216 560654 510258 566772
rect 510494 560654 510536 566772
rect 512421 566697 515308 567251
rect 517160 567176 517202 573294
rect 517438 567176 517480 573294
rect 519350 573219 522237 573773
rect 517800 573195 523768 573219
rect 517800 567275 517824 573195
rect 519350 567275 522237 573195
rect 523744 567275 523768 573195
rect 517800 567251 523768 567275
rect 517160 566772 517480 567176
rect 510856 566673 516824 566697
rect 510856 560753 510880 566673
rect 512421 560753 515308 566673
rect 516800 560753 516824 566673
rect 510856 560729 516824 560753
rect 510216 560452 510536 560654
rect 512421 555373 515308 560729
rect 517160 560654 517202 566772
rect 517438 560654 517480 566772
rect 519350 566697 522237 567251
rect 517800 566673 523768 566697
rect 517800 560753 517824 566673
rect 519350 560753 522237 566673
rect 523744 560753 523768 566673
rect 517800 560729 523768 560753
rect 517160 560452 517480 560654
rect 519350 555373 522237 560729
rect 491289 555225 522237 555373
rect 491289 540589 491316 555225
rect 521952 540589 522237 555225
rect 491289 540442 522237 540589
rect 451976 378829 467642 540237
rect 519350 540149 522237 540442
rect 451976 363553 452175 378829
rect 467131 363553 467642 378829
rect 451976 240343 467642 363553
rect 451976 227015 452145 240343
rect 452007 225387 452145 227015
rect 467421 227015 467642 240343
rect 545384 432002 561540 584115
rect 545384 417366 545733 432002
rect 561009 417366 561540 432002
rect 467421 225387 467559 227015
rect 452007 225352 467559 225387
rect 338385 136722 338714 151535
rect 100463 136311 116619 136634
rect 338617 136579 338714 136722
rect 354310 136722 354541 151535
rect 545384 151638 561540 417366
rect 545384 137728 545507 151638
rect 354310 136579 354407 136722
rect 545458 136682 545507 137728
rect 561423 137728 561540 151638
rect 561423 136682 561472 137728
rect 545458 136595 561472 136682
rect 338617 136437 354407 136579
use mimcap_decoup_1x5  mimcap_decoup_1x5_6
array 0 0 34500 0 2 6522
timestamp 1624397418
transform 1 0 38481 0 1 560871
box 0 -159 34500 6363
use top_pll_v1  top_pll_v1_1
timestamp 1624397418
transform 1 0 14782 0 1 657248
box -656 -33693 50195 2860
use sky130_fd_pr__cap_mim_m3_2_2Y8F6P  sky130_fd_pr__cap_mim_m3_2_2Y8F6P_2
array 0 0 6724 0 8 6522
timestamp 1624397418
transform 1 0 74005 0 1 616157
box -3351 -3261 3373 3261
use top_pll_v2  top_pll_v2_0
timestamp 1624397418
transform -1 0 133068 0 1 657248
box -656 -33693 50195 2860
use mimcap_decoup_1x5  mimcap_decoup_1x5_5
array 0 0 34500 0 2 6522
timestamp 1624397418
transform 1 0 126717 0 1 559996
box 0 -159 34500 6363
use sky130_fd_pr__cap_mim_m3_2_2Y8F6P  sky130_fd_pr__cap_mim_m3_2_2Y8F6P_1
array 0 0 6724 0 8 6522
timestamp 1624397418
transform 1 0 144463 0 1 616442
box -3351 -3261 3373 3261
use top_pll_v1  top_pll_v1_0
timestamp 1624397418
transform -1 0 206380 0 1 656706
box -656 -33693 50195 2860
use sky130_fd_pr__cap_mim_m3_2_2Y8F6P  sky130_fd_pr__cap_mim_m3_2_2Y8F6P_0
array 0 0 6724 0 6 6522
timestamp 1624397418
transform 1 0 220679 0 1 616773
box -3351 -3261 3373 3261
use mimcap_decoup_1x5  mimcap_decoup_1x5_4
array 0 0 34500 0 2 6522
timestamp 1624397418
transform 1 0 197202 0 1 560156
box 0 -159 34500 6363
use bias  bias_0
timestamp 1624397418
transform 1 0 202834 0 -1 687483
box -54 -412 44317 2238
use mimcap_decoup_1x5  mimcap_decoup_1x5_3
array 0 0 34500 0 1 6522
timestamp 1624397418
transform -1 0 345445 0 1 602155
box 0 -159 34500 6363
use mimcap_decoup_1x5  mimcap_decoup_1x5_2
array 0 0 34500 0 2 6522
timestamp 1624397418
transform 1 0 291410 0 1 559700
box 0 -159 34500 6363
use res_amp_top  res_amp_top_0
timestamp 1624397418
transform 1 0 349695 0 1 630386
box -5005 -972 31038 12726
use mimcap_decoup_1x5  mimcap_decoup_1x5_1
array 0 0 34500 0 2 6522
timestamp 1624397418
transform 1 0 382888 0 1 560156
box 0 -159 34500 6363
use mimcap_decoup_1x5  mimcap_decoup_1x5_0
array 0 0 34500 0 2 6522
timestamp 1624397418
transform 1 0 489384 0 1 560611
box 0 -159 34500 6363
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s -800 559442 860 564242 0 FreeSans 1400 180 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
