magic
tech sky130A
magscale 1 2
timestamp 1624065706
<< nwell >>
rect -422 2867 0 2956
<< pwell >>
rect 1294 809 1725 1389
rect 2588 809 3019 1389
rect -422 165 -411 166
rect -422 0 0 165
<< psubdiff >>
rect -314 36 -290 70
rect -132 36 -108 70
<< nsubdiff >>
rect -314 2886 -290 2920
rect -132 2886 -108 2920
<< psubdiffcont >>
rect -290 36 -132 70
<< nsubdiffcont >>
rect -290 2886 -132 2920
<< viali >>
rect -386 2886 -290 2920
rect -290 2886 -132 2920
rect -132 2886 -36 2920
rect -386 2797 -36 2831
rect -386 125 -36 159
rect -386 36 -290 70
rect -290 36 -132 70
rect -132 36 -36 70
<< metal1 >>
rect -422 2920 3882 2926
rect -422 2886 -386 2920
rect -36 2898 3882 2920
rect -36 2886 0 2898
rect -422 2831 0 2886
rect -422 2797 -386 2831
rect -36 2797 0 2831
rect -422 2791 0 2797
rect -324 2348 -278 2791
rect -243 2695 -233 2747
rect -129 2695 -119 2747
rect 1264 2738 1323 2781
rect 2559 2738 2625 2801
rect 3873 2738 3882 2778
rect -243 2686 -144 2695
rect -190 2646 -144 2686
rect -190 2199 -144 2353
rect -236 739 -98 2199
rect 1294 783 1725 957
rect 2588 783 3019 957
rect 1294 779 1727 783
rect 2588 779 3021 783
rect 1295 746 1727 779
rect 2589 746 3021 779
rect -324 165 -278 599
rect -190 597 -144 739
rect -243 261 -119 270
rect -243 209 -233 261
rect -129 209 -119 261
rect -422 159 0 165
rect -422 125 -386 159
rect -36 125 0 159
rect -422 70 0 125
rect 686 70 3266 165
rect -422 36 -386 70
rect -36 36 0 70
rect -422 30 0 36
<< via1 >>
rect -233 2695 -129 2747
rect -233 209 -129 261
<< metal2 >>
rect -233 2747 3266 2757
rect -129 2695 3266 2747
rect -233 2685 3266 2695
rect 443 2631 678 2685
rect 1736 2631 1971 2685
rect 3031 2638 3266 2685
rect 440 1417 608 1427
rect 3316 1417 3440 1427
rect 1255 1363 1757 1415
rect 2557 1363 3030 1415
rect 440 1351 608 1361
rect 3651 1363 3882 1415
rect 3316 1351 3440 1361
rect 436 299 678 300
rect 436 278 684 299
rect -230 271 684 278
rect -233 261 684 271
rect -129 209 684 261
rect -233 199 684 209
rect -230 184 684 199
rect 564 162 684 184
rect 1730 162 1971 295
rect 3023 162 3214 294
rect 564 68 3215 162
<< via2 >>
rect 440 1361 608 1417
rect 3316 1361 3440 1417
<< metal3 >>
rect 430 1421 618 1422
rect 430 1417 441 1421
rect 607 1417 618 1421
rect 430 1361 440 1417
rect 608 1361 618 1417
rect 430 1357 441 1361
rect 607 1357 618 1361
rect 430 1356 618 1357
rect 3306 1421 3450 1425
rect 3306 1417 3317 1421
rect 3306 1361 3316 1417
rect 3306 1357 3317 1361
rect 3440 1357 3450 1421
rect 3306 1353 3450 1357
rect 3601 868 3661 1007
rect 983 797 993 868
rect 1100 797 1110 868
rect 2289 799 2299 867
rect 2377 799 2387 867
rect 3584 799 3594 866
rect 3672 799 3682 866
rect 3601 88 3661 799
<< via3 >>
rect 441 1417 607 1421
rect 441 1361 607 1417
rect 441 1357 607 1361
rect 3317 1417 3440 1421
rect 3317 1361 3440 1417
rect 3317 1357 3440 1361
rect 993 797 1100 868
rect 2299 799 2377 867
rect 3594 799 3672 866
<< metal4 >>
rect 440 1421 608 1422
rect 3316 1421 3441 1422
rect 440 1357 441 1421
rect 607 1357 3317 1421
rect 3440 1357 3441 1421
rect 440 1356 608 1357
rect 3316 1356 3441 1357
rect 992 868 3680 869
rect 992 797 993 868
rect 1100 867 3680 868
rect 1100 799 2299 867
rect 2377 866 3680 867
rect 2377 799 3594 866
rect 3672 799 3680 866
rect 1100 798 3680 799
rect 1100 797 1101 798
rect 992 796 1101 797
use csvco_branch_v2  csvco_branch_v2_1
timestamp 1624064496
transform 1 0 1657 0 1 1002
box -363 -1002 932 1955
use csvco_branch_v2  csvco_branch_v2_2
timestamp 1624064496
transform 1 0 2951 0 1 1002
box -363 -1002 932 1955
use sky130_fd_pr__pfet_01v8_4757AC  sky130_fd_pr__pfet_01v8_4757AC_0
timestamp 1624049879
transform 1 0 -211 0 1 2498
box -211 -369 211 369
use sky130_fd_pr__nfet_01v8_CBAU6Y  sky130_fd_pr__nfet_01v8_CBAU6Y_0
timestamp 1624049879
transform 1 0 -211 0 1 449
box -211 -360 211 360
use csvco_branch_v2  csvco_branch_v2_0
timestamp 1624064496
transform 1 0 363 0 1 1002
box -363 -1002 932 1955
<< labels >>
rlabel metal1 -422 70 0 125 1 vss
rlabel metal1 -422 2831 0 2886 1 vdd
rlabel metal2 3651 1363 3882 1415 1 out_vco
rlabel metal3 3601 88 3661 148 1 D0
rlabel metal2 -105 212 -39 260 1 vctrl
rlabel metal2 41 2699 69 2726 1 vbp
<< end >>
