magic
tech sky130A
magscale 1 2
timestamp 1624043228
<< pwell >>
rect 2250 1287 5928 1291
rect 2049 850 2193 1059
rect 2250 621 5928 625
rect 2250 355 5928 359
rect 2250 -1147 5928 -1143
rect 6242 -1261 6276 1390
rect 7186 -616 7209 -612
rect 372 -1391 2014 -1357
rect 2086 -1392 6188 -1358
<< psubdiff >>
rect 6242 1343 6276 1390
rect 6242 411 6276 569
rect 6242 -1261 6276 -1199
rect 372 -1391 468 -1357
rect 1114 -1391 1272 -1357
rect 1918 -1391 2014 -1357
rect 2086 -1392 2182 -1358
rect 6092 -1392 6188 -1358
<< psubdiffcont >>
rect 6242 569 6276 1343
rect 6242 -1199 6276 411
rect 468 -1391 1114 -1357
rect 1272 -1391 1918 -1357
rect 2182 -1392 6092 -1358
<< poly >>
rect 2250 1287 2280 1291
rect 2346 1287 2376 1291
rect 2442 1287 2472 1291
rect 2538 1287 2568 1291
rect 2634 1287 2664 1291
rect 2730 1287 2760 1291
rect 2826 1287 2856 1291
rect 2922 1287 2952 1291
rect 3018 1287 3048 1291
rect 3114 1287 3144 1291
rect 3210 1287 3240 1291
rect 3306 1287 3336 1291
rect 3402 1287 3432 1291
rect 3498 1287 3528 1291
rect 3594 1287 3624 1291
rect 3690 1287 3720 1291
rect 3786 1287 3816 1291
rect 3882 1287 3912 1291
rect 3978 1287 4008 1291
rect 4074 1287 4104 1291
rect 4170 1287 4200 1291
rect 4266 1287 4296 1291
rect 4362 1287 4392 1291
rect 4458 1287 4488 1291
rect 4554 1287 4584 1291
rect 4650 1287 4680 1291
rect 4746 1287 4776 1291
rect 4842 1287 4872 1291
rect 4938 1287 4968 1291
rect 5034 1287 5064 1291
rect 5130 1287 5160 1291
rect 5226 1287 5256 1291
rect 5322 1287 5352 1291
rect 5418 1287 5448 1291
rect 5514 1287 5544 1291
rect 5610 1287 5640 1291
rect 5706 1287 5736 1291
rect 5802 1287 5832 1291
rect 5898 1287 5928 1291
rect 2068 1024 2235 1043
rect 2068 890 2083 1024
rect 2129 890 2235 1024
rect 2068 869 2235 890
rect 2250 621 2280 625
rect 2346 621 2376 625
rect 2442 621 2472 625
rect 2538 621 2568 625
rect 2634 621 2664 625
rect 2730 621 2760 625
rect 2826 621 2856 625
rect 2922 621 2952 625
rect 3018 621 3048 625
rect 3114 621 3144 625
rect 3210 621 3240 625
rect 3306 621 3336 625
rect 3402 621 3432 625
rect 3498 621 3528 625
rect 3594 621 3624 625
rect 3690 621 3720 625
rect 3786 621 3816 625
rect 3882 621 3912 625
rect 3978 621 4008 625
rect 4074 621 4104 625
rect 4170 621 4200 625
rect 4266 621 4296 625
rect 4362 621 4392 625
rect 4458 621 4488 625
rect 4554 621 4584 625
rect 4650 621 4680 625
rect 4746 621 4776 625
rect 4842 621 4872 625
rect 4938 621 4968 625
rect 5034 621 5064 625
rect 5130 621 5160 625
rect 5226 621 5256 625
rect 5322 621 5352 625
rect 5418 621 5448 625
rect 5514 621 5544 625
rect 5610 621 5640 625
rect 5706 621 5736 625
rect 5802 621 5832 625
rect 5898 621 5928 625
rect 2250 355 2280 359
rect 2346 355 2376 359
rect 2442 355 2472 359
rect 2538 355 2568 359
rect 2634 355 2664 359
rect 2730 355 2760 359
rect 2826 355 2856 359
rect 2922 355 2952 359
rect 3018 355 3048 359
rect 3114 355 3144 359
rect 3210 355 3240 359
rect 3306 355 3336 359
rect 3402 355 3432 359
rect 3498 355 3528 359
rect 3594 355 3624 359
rect 3690 355 3720 359
rect 3786 355 3816 359
rect 3882 355 3912 359
rect 3978 355 4008 359
rect 4074 355 4104 359
rect 4170 355 4200 359
rect 4266 355 4296 359
rect 4362 355 4392 359
rect 4458 355 4488 359
rect 4554 355 4584 359
rect 4650 355 4680 359
rect 4746 355 4776 359
rect 4842 355 4872 359
rect 4938 355 4968 359
rect 5034 355 5064 359
rect 5130 355 5160 359
rect 5226 355 5256 359
rect 5322 355 5352 359
rect 5418 355 5448 359
rect 5514 355 5544 359
rect 5610 355 5640 359
rect 5706 355 5736 359
rect 5802 355 5832 359
rect 5898 355 5928 359
rect 2069 92 2259 111
rect 2069 -42 2084 92
rect 2130 -42 2259 92
rect 2069 -63 2259 -42
rect 2069 -326 2259 -307
rect 2069 -460 2084 -326
rect 2130 -460 2259 -326
rect 2069 -481 2259 -460
rect 2069 -744 2259 -725
rect 2069 -878 2084 -744
rect 2130 -878 2259 -744
rect 2069 -899 2259 -878
rect 2250 -1147 2280 -1143
rect 2346 -1147 2376 -1143
rect 2442 -1147 2472 -1143
rect 2538 -1147 2568 -1143
rect 2634 -1147 2664 -1143
rect 2730 -1147 2760 -1143
rect 2826 -1147 2856 -1143
rect 2922 -1147 2952 -1143
rect 3018 -1147 3048 -1143
rect 3114 -1147 3144 -1143
rect 3210 -1147 3240 -1143
rect 3306 -1147 3336 -1143
rect 3402 -1147 3432 -1143
rect 3498 -1147 3528 -1143
rect 3594 -1147 3624 -1143
rect 3690 -1147 3720 -1143
rect 3786 -1147 3816 -1143
rect 3882 -1147 3912 -1143
rect 3978 -1147 4008 -1143
rect 4074 -1147 4104 -1143
rect 4170 -1147 4200 -1143
rect 4266 -1147 4296 -1143
rect 4362 -1147 4392 -1143
rect 4458 -1147 4488 -1143
rect 4554 -1147 4584 -1143
rect 4650 -1147 4680 -1143
rect 4746 -1147 4776 -1143
rect 4842 -1147 4872 -1143
rect 4938 -1147 4968 -1143
rect 5034 -1147 5064 -1143
rect 5130 -1147 5160 -1143
rect 5226 -1147 5256 -1143
rect 5322 -1147 5352 -1143
rect 5418 -1147 5448 -1143
rect 5514 -1147 5544 -1143
rect 5610 -1147 5640 -1143
rect 5706 -1147 5736 -1143
rect 5802 -1147 5832 -1143
rect 5898 -1147 5928 -1143
<< polycont >>
rect 2083 890 2129 1024
rect 2084 -42 2130 92
rect 2084 -460 2130 -326
rect 2084 -878 2130 -744
<< viali >>
rect 2083 1024 2129 1043
rect 2083 890 2129 1024
rect 2083 869 2129 890
rect 2084 92 2130 111
rect 2084 -42 2130 92
rect 2084 -63 2130 -42
rect 2084 -326 2130 -307
rect 2084 -460 2130 -326
rect 2084 -481 2130 -460
rect 2084 -744 2130 -725
rect 2084 -878 2130 -744
rect 2084 -899 2130 -878
rect 6154 -1261 6188 1390
rect 6242 1343 6276 1390
rect 6242 569 6276 1343
rect 6242 411 6276 569
rect 6242 -1199 6276 411
rect 6242 -1261 6276 -1199
rect 372 -1303 2014 -1269
rect 2086 -1295 6188 -1261
rect 372 -1391 468 -1357
rect 468 -1391 1114 -1357
rect 1114 -1391 1272 -1357
rect 1272 -1391 1918 -1357
rect 1918 -1391 2014 -1357
rect 2086 -1392 2182 -1358
rect 2182 -1392 6092 -1358
rect 6092 -1392 6188 -1358
<< metal1 >>
rect 2194 1405 6080 1545
rect 2010 1043 2135 1055
rect 2010 869 2083 1043
rect 2129 869 2135 1043
rect 2010 850 2135 869
rect 2194 647 2240 1405
rect 2270 1065 2280 1265
rect 2346 1065 2356 1265
rect 2270 647 2280 847
rect 2346 647 2356 847
rect 2386 647 2432 1405
rect 2462 1065 2472 1265
rect 2538 1065 2548 1265
rect 2462 647 2472 847
rect 2538 647 2548 847
rect 2578 647 2624 1405
rect 2654 1065 2664 1265
rect 2730 1065 2740 1265
rect 2654 647 2664 847
rect 2730 647 2740 847
rect 2770 647 2816 1405
rect 2846 1065 2856 1265
rect 2922 1065 2932 1265
rect 2846 647 2856 847
rect 2922 647 2932 847
rect 2962 647 3008 1405
rect 3038 1065 3048 1265
rect 3114 1065 3124 1265
rect 3038 647 3048 847
rect 3114 647 3124 847
rect 3154 647 3200 1405
rect 3230 1065 3240 1265
rect 3306 1065 3316 1265
rect 3230 647 3240 847
rect 3306 647 3316 847
rect 3346 647 3392 1405
rect 3422 1065 3432 1265
rect 3498 1065 3508 1265
rect 3422 647 3432 847
rect 3498 647 3508 847
rect 3538 647 3584 1405
rect 3614 1065 3624 1265
rect 3690 1065 3700 1265
rect 3614 647 3624 847
rect 3690 647 3700 847
rect 3730 647 3776 1405
rect 3806 1065 3816 1265
rect 3882 1065 3892 1265
rect 3806 647 3816 847
rect 3882 647 3892 847
rect 3922 647 3968 1405
rect 3998 1065 4008 1265
rect 4074 1065 4084 1265
rect 3998 647 4008 847
rect 4074 647 4084 847
rect 4114 647 4160 1405
rect 4190 1065 4200 1265
rect 4266 1065 4276 1265
rect 4190 647 4200 847
rect 4266 647 4276 847
rect 4306 647 4352 1405
rect 4382 1065 4392 1265
rect 4458 1065 4468 1265
rect 4382 647 4392 847
rect 4458 647 4468 847
rect 4498 647 4544 1405
rect 4574 1065 4584 1265
rect 4650 1065 4660 1265
rect 4574 647 4584 847
rect 4650 647 4660 847
rect 4690 647 4736 1405
rect 4766 1065 4776 1265
rect 4842 1065 4852 1265
rect 4766 647 4776 847
rect 4842 647 4852 847
rect 4882 647 4928 1405
rect 4958 1065 4968 1265
rect 5034 1065 5044 1265
rect 4958 647 4968 847
rect 5034 647 5044 847
rect 5074 647 5120 1405
rect 5150 1065 5160 1265
rect 5226 1065 5236 1265
rect 5150 647 5160 847
rect 5226 647 5236 847
rect 5266 647 5312 1405
rect 5342 1065 5352 1265
rect 5418 1065 5428 1265
rect 5342 647 5352 847
rect 5418 647 5428 847
rect 5458 647 5504 1405
rect 5534 1065 5544 1265
rect 5610 1065 5620 1265
rect 5534 647 5544 847
rect 5610 647 5620 847
rect 5650 647 5696 1405
rect 5726 1065 5736 1265
rect 5802 1065 5812 1265
rect 5726 647 5736 847
rect 5802 647 5812 847
rect 5842 647 5888 1405
rect 5918 1065 5928 1265
rect 5994 1065 6004 1265
rect 5918 647 5928 847
rect 5994 647 6004 847
rect 6034 647 6080 1405
rect 6147 1390 6282 1402
rect 2069 111 2136 123
rect 1961 -63 2084 111
rect 2130 -63 2136 111
rect 1961 -307 2136 -63
rect 1961 -481 2084 -307
rect 2130 -481 2136 -307
rect 1961 -713 2136 -481
rect 520 -725 2136 -713
rect 520 -899 2084 -725
rect 2130 -899 2136 -725
rect 520 -901 2136 -899
rect 460 -1129 470 -929
rect 536 -1129 546 -929
rect 576 -933 622 -901
rect 652 -1129 662 -929
rect 728 -1129 738 -929
rect 768 -933 814 -901
rect 844 -1129 854 -929
rect 920 -1129 930 -929
rect 960 -939 1006 -901
rect 2069 -911 2136 -901
rect 1036 -1129 1046 -929
rect 1112 -1129 1122 -929
rect 1284 -1253 1330 -1105
rect 1360 -1129 1370 -929
rect 1436 -1129 1446 -929
rect 1476 -1253 1522 -1102
rect 1552 -1129 1562 -929
rect 1628 -1129 1638 -929
rect 1668 -1253 1714 -1108
rect 1744 -1129 1754 -929
rect 1820 -1129 1830 -929
rect 1860 -1253 1906 -1116
rect 2194 -1253 2240 291
rect 2270 133 2280 333
rect 2346 133 2356 333
rect 2270 -285 2280 -85
rect 2346 -285 2356 -85
rect 2270 -703 2280 -503
rect 2346 -703 2356 -503
rect 2270 -1121 2280 -921
rect 2346 -1121 2356 -921
rect 2386 -1253 2432 299
rect 2462 133 2472 333
rect 2538 133 2548 333
rect 2462 -285 2472 -85
rect 2538 -285 2548 -85
rect 2462 -703 2472 -503
rect 2538 -703 2548 -503
rect 2462 -1121 2472 -921
rect 2538 -1121 2548 -921
rect 2578 -1253 2624 297
rect 2654 133 2664 333
rect 2730 133 2740 333
rect 2654 -285 2664 -85
rect 2730 -285 2740 -85
rect 2654 -703 2664 -503
rect 2730 -703 2740 -503
rect 2654 -1121 2664 -921
rect 2730 -1121 2740 -921
rect 2770 -1253 2816 301
rect 2846 133 2856 333
rect 2922 133 2932 333
rect 2846 -285 2856 -85
rect 2922 -285 2932 -85
rect 2846 -703 2856 -503
rect 2922 -703 2932 -503
rect 2846 -1121 2856 -921
rect 2922 -1121 2932 -921
rect 2962 -1253 3008 270
rect 3038 133 3048 333
rect 3114 133 3124 333
rect 3038 -285 3048 -85
rect 3114 -285 3124 -85
rect 3038 -703 3048 -503
rect 3114 -703 3124 -503
rect 3038 -1121 3048 -921
rect 3114 -1121 3124 -921
rect 3154 -1253 3200 278
rect 3230 133 3240 333
rect 3306 133 3316 333
rect 3230 -285 3240 -85
rect 3306 -285 3316 -85
rect 3230 -703 3240 -503
rect 3306 -703 3316 -503
rect 3230 -1121 3240 -921
rect 3306 -1121 3316 -921
rect 3346 -1253 3392 277
rect 3422 133 3432 333
rect 3498 133 3508 333
rect 3422 -285 3432 -85
rect 3498 -285 3508 -85
rect 3422 -703 3432 -503
rect 3498 -703 3508 -503
rect 3422 -1121 3432 -921
rect 3498 -1121 3508 -921
rect 3539 -1253 3585 279
rect 3614 133 3624 333
rect 3690 133 3700 333
rect 3614 -285 3624 -85
rect 3690 -285 3700 -85
rect 3614 -703 3624 -503
rect 3690 -703 3700 -503
rect 3614 -1121 3624 -921
rect 3690 -1121 3700 -921
rect 3730 -1253 3776 273
rect 3806 133 3816 333
rect 3882 133 3892 333
rect 3806 -285 3816 -85
rect 3882 -285 3892 -85
rect 3806 -703 3816 -503
rect 3882 -703 3892 -503
rect 3806 -1121 3816 -921
rect 3882 -1121 3892 -921
rect 3922 -1253 3968 281
rect 3998 133 4008 333
rect 4074 133 4084 333
rect 3998 -285 4008 -85
rect 4074 -285 4084 -85
rect 3998 -703 4008 -503
rect 4074 -703 4084 -503
rect 3998 -1121 4008 -921
rect 4074 -1121 4084 -921
rect 4114 -1253 4160 282
rect 4190 133 4200 333
rect 4266 133 4276 333
rect 4190 -285 4200 -85
rect 4266 -285 4276 -85
rect 4190 -703 4200 -503
rect 4266 -703 4276 -503
rect 4190 -1121 4200 -921
rect 4266 -1121 4276 -921
rect 4306 -1253 4352 281
rect 4382 133 4392 333
rect 4458 133 4468 333
rect 4382 -285 4392 -85
rect 4458 -285 4468 -85
rect 4382 -703 4392 -503
rect 4458 -703 4468 -503
rect 4382 -1121 4392 -921
rect 4458 -1121 4468 -921
rect 4498 -1253 4544 282
rect 4574 133 4584 333
rect 4650 133 4660 333
rect 4574 -285 4584 -85
rect 4650 -285 4660 -85
rect 4574 -703 4584 -503
rect 4650 -703 4660 -503
rect 4574 -1121 4584 -921
rect 4650 -1121 4660 -921
rect 4690 -1253 4736 280
rect 4766 133 4776 333
rect 4842 133 4852 333
rect 4766 -285 4776 -85
rect 4842 -285 4852 -85
rect 4766 -703 4776 -503
rect 4842 -703 4852 -503
rect 4766 -1121 4776 -921
rect 4842 -1121 4852 -921
rect 4882 -1253 4928 279
rect 4958 133 4968 333
rect 5034 133 5044 333
rect 4958 -285 4968 -85
rect 5034 -285 5044 -85
rect 4958 -703 4968 -503
rect 5034 -703 5044 -503
rect 4958 -1121 4968 -921
rect 5034 -1121 5044 -921
rect 5074 -1253 5120 277
rect 5150 133 5160 333
rect 5226 133 5236 333
rect 5150 -285 5160 -85
rect 5226 -285 5236 -85
rect 5150 -703 5160 -503
rect 5226 -703 5236 -503
rect 5150 -1121 5160 -921
rect 5226 -1121 5236 -921
rect 5266 -1253 5312 277
rect 5342 133 5352 333
rect 5418 133 5428 333
rect 5342 -285 5352 -85
rect 5418 -285 5428 -85
rect 5342 -703 5352 -503
rect 5418 -703 5428 -503
rect 5342 -1121 5352 -921
rect 5418 -1121 5428 -921
rect 5458 -1253 5504 279
rect 5534 133 5544 333
rect 5610 133 5620 333
rect 5534 -285 5544 -85
rect 5610 -285 5620 -85
rect 5534 -703 5544 -503
rect 5610 -703 5620 -503
rect 5534 -1121 5544 -921
rect 5610 -1121 5620 -921
rect 5650 -1253 5696 275
rect 5726 133 5736 333
rect 5802 133 5812 333
rect 5726 -285 5736 -85
rect 5802 -285 5812 -85
rect 5726 -703 5736 -503
rect 5802 -703 5812 -503
rect 5726 -1121 5736 -921
rect 5802 -1121 5812 -921
rect 5842 -1253 5888 277
rect 5918 133 5928 333
rect 5994 133 6004 333
rect 5918 -285 5928 -85
rect 5994 -285 6004 -85
rect 5918 -703 5928 -503
rect 5994 -703 6004 -503
rect 5918 -1121 5928 -921
rect 5994 -1121 6004 -921
rect 6034 -1253 6080 274
rect 6147 -1253 6154 1390
rect 336 -1261 6154 -1253
rect 6188 -1261 6242 1390
rect 6276 -1261 6282 1390
rect 336 -1269 2086 -1261
rect 336 -1303 372 -1269
rect 2014 -1295 2086 -1269
rect 6188 -1295 6282 -1261
rect 2014 -1303 6282 -1295
rect 336 -1357 6282 -1303
rect 336 -1391 372 -1357
rect 2014 -1358 6282 -1357
rect 2014 -1391 2086 -1358
rect 336 -1392 2086 -1391
rect 6188 -1392 6282 -1358
rect 336 -1409 6282 -1392
<< via1 >>
rect 2280 1065 2346 1265
rect 2280 647 2346 847
rect 2472 1065 2538 1265
rect 2472 647 2538 847
rect 2664 1065 2730 1265
rect 2664 647 2730 847
rect 2856 1065 2922 1265
rect 2856 647 2922 847
rect 3048 1065 3114 1265
rect 3048 647 3114 847
rect 3240 1065 3306 1265
rect 3240 647 3306 847
rect 3432 1065 3498 1265
rect 3432 647 3498 847
rect 3624 1065 3690 1265
rect 3624 647 3690 847
rect 3816 1065 3882 1265
rect 3816 647 3882 847
rect 4008 1065 4074 1265
rect 4008 647 4074 847
rect 4200 1065 4266 1265
rect 4200 647 4266 847
rect 4392 1065 4458 1265
rect 4392 647 4458 847
rect 4584 1065 4650 1265
rect 4584 647 4650 847
rect 4776 1065 4842 1265
rect 4776 647 4842 847
rect 4968 1065 5034 1265
rect 4968 647 5034 847
rect 5160 1065 5226 1265
rect 5160 647 5226 847
rect 5352 1065 5418 1265
rect 5352 647 5418 847
rect 5544 1065 5610 1265
rect 5544 647 5610 847
rect 5736 1065 5802 1265
rect 5736 647 5802 847
rect 5928 1065 5994 1265
rect 5928 647 5994 847
rect 470 -1129 536 -929
rect 662 -1129 728 -929
rect 854 -1129 920 -929
rect 1046 -1129 1112 -929
rect 1370 -1129 1436 -929
rect 1562 -1129 1628 -929
rect 1754 -1129 1820 -929
rect 2280 133 2346 333
rect 2280 -285 2346 -85
rect 2280 -703 2346 -503
rect 2280 -1121 2346 -921
rect 2472 133 2538 333
rect 2472 -285 2538 -85
rect 2472 -703 2538 -503
rect 2472 -1121 2538 -921
rect 2664 133 2730 333
rect 2664 -285 2730 -85
rect 2664 -703 2730 -503
rect 2664 -1121 2730 -921
rect 2856 133 2922 333
rect 2856 -285 2922 -85
rect 2856 -703 2922 -503
rect 2856 -1121 2922 -921
rect 3048 133 3114 333
rect 3048 -285 3114 -85
rect 3048 -703 3114 -503
rect 3048 -1121 3114 -921
rect 3240 133 3306 333
rect 3240 -285 3306 -85
rect 3240 -703 3306 -503
rect 3240 -1121 3306 -921
rect 3432 133 3498 333
rect 3432 -285 3498 -85
rect 3432 -703 3498 -503
rect 3432 -1121 3498 -921
rect 3624 133 3690 333
rect 3624 -285 3690 -85
rect 3624 -703 3690 -503
rect 3624 -1121 3690 -921
rect 3816 133 3882 333
rect 3816 -285 3882 -85
rect 3816 -703 3882 -503
rect 3816 -1121 3882 -921
rect 4008 133 4074 333
rect 4008 -285 4074 -85
rect 4008 -703 4074 -503
rect 4008 -1121 4074 -921
rect 4200 133 4266 333
rect 4200 -285 4266 -85
rect 4200 -703 4266 -503
rect 4200 -1121 4266 -921
rect 4392 133 4458 333
rect 4392 -285 4458 -85
rect 4392 -703 4458 -503
rect 4392 -1121 4458 -921
rect 4584 133 4650 333
rect 4584 -285 4650 -85
rect 4584 -703 4650 -503
rect 4584 -1121 4650 -921
rect 4776 133 4842 333
rect 4776 -285 4842 -85
rect 4776 -703 4842 -503
rect 4776 -1121 4842 -921
rect 4968 133 5034 333
rect 4968 -285 5034 -85
rect 4968 -703 5034 -503
rect 4968 -1121 5034 -921
rect 5160 133 5226 333
rect 5160 -285 5226 -85
rect 5160 -703 5226 -503
rect 5160 -1121 5226 -921
rect 5352 133 5418 333
rect 5352 -285 5418 -85
rect 5352 -703 5418 -503
rect 5352 -1121 5418 -921
rect 5544 133 5610 333
rect 5544 -285 5610 -85
rect 5544 -703 5610 -503
rect 5544 -1121 5610 -921
rect 5736 133 5802 333
rect 5736 -285 5802 -85
rect 5736 -703 5802 -503
rect 5736 -1121 5802 -921
rect 5928 133 5994 333
rect 5928 -285 5994 -85
rect 5928 -703 5994 -503
rect 5928 -1121 5994 -921
<< metal2 >>
rect 2280 1265 2346 1275
rect 2280 847 2346 1065
rect 2280 596 2346 647
rect 2472 1265 2538 1275
rect 2472 847 2538 1065
rect 2472 596 2538 647
rect 2664 1265 2730 1275
rect 2664 847 2730 1065
rect 2664 596 2730 647
rect 2856 1265 2922 1275
rect 2856 847 2922 1065
rect 2856 596 2922 647
rect 3048 1265 3114 1275
rect 3048 847 3114 1065
rect 3048 596 3114 647
rect 3240 1265 3306 1275
rect 3240 847 3306 1065
rect 3240 596 3306 647
rect 3432 1265 3498 1275
rect 3432 847 3498 1065
rect 3432 596 3498 647
rect 3624 1265 3690 1275
rect 3624 847 3690 1065
rect 3624 596 3690 647
rect 3816 1265 3882 1275
rect 3816 847 3882 1065
rect 3816 596 3882 647
rect 4008 1265 4074 1275
rect 4008 847 4074 1065
rect 4008 596 4074 647
rect 4200 1265 4266 1275
rect 4200 847 4266 1065
rect 4200 596 4266 647
rect 4392 1265 4458 1275
rect 4392 847 4458 1065
rect 4392 596 4458 647
rect 4584 1265 4650 1275
rect 4584 847 4650 1065
rect 4584 596 4650 647
rect 4776 1265 4842 1275
rect 4776 847 4842 1065
rect 4776 596 4842 647
rect 4968 1265 5034 1275
rect 4968 847 5034 1065
rect 4968 596 5034 647
rect 5160 1265 5226 1275
rect 5160 847 5226 1065
rect 5160 596 5226 647
rect 5352 1265 5418 1275
rect 5352 847 5418 1065
rect 5352 596 5418 647
rect 5544 1265 5610 1275
rect 5544 847 5610 1065
rect 5544 596 5610 647
rect 5736 1265 5802 1275
rect 5736 847 5802 1065
rect 5736 596 5802 647
rect 5928 1265 5994 1275
rect 5928 847 5994 1065
rect 5928 596 5994 647
rect 2280 389 5994 596
rect 2280 333 2346 389
rect 2280 -85 2346 133
rect 2280 -503 2346 -285
rect 470 -929 1820 -919
rect 536 -1129 662 -929
rect 728 -1129 854 -929
rect 920 -1129 1046 -929
rect 1112 -1129 1370 -929
rect 1436 -1129 1562 -929
rect 1628 -1129 1754 -929
rect 470 -1139 1820 -1129
rect 2280 -921 2346 -703
rect 2280 -1131 2346 -1121
rect 2472 333 2538 389
rect 2472 -85 2538 133
rect 2472 -503 2538 -285
rect 2472 -921 2538 -703
rect 2472 -1131 2538 -1121
rect 2664 333 2730 389
rect 2664 -85 2730 133
rect 2664 -503 2730 -285
rect 2664 -921 2730 -703
rect 2664 -1131 2730 -1121
rect 2856 333 2922 389
rect 2856 -85 2922 133
rect 2856 -503 2922 -285
rect 2856 -921 2922 -703
rect 2856 -1131 2922 -1121
rect 3048 333 3114 389
rect 3048 -85 3114 133
rect 3048 -503 3114 -285
rect 3048 -921 3114 -703
rect 3048 -1131 3114 -1121
rect 3240 333 3306 389
rect 3240 -85 3306 133
rect 3240 -503 3306 -285
rect 3240 -921 3306 -703
rect 3240 -1131 3306 -1121
rect 3432 333 3498 389
rect 3432 -85 3498 133
rect 3432 -503 3498 -285
rect 3432 -921 3498 -703
rect 3432 -1131 3498 -1121
rect 3624 333 3690 389
rect 3624 -85 3690 133
rect 3624 -503 3690 -285
rect 3624 -921 3690 -703
rect 3624 -1131 3690 -1121
rect 3816 333 3882 389
rect 3816 -85 3882 133
rect 3816 -503 3882 -285
rect 3816 -921 3882 -703
rect 3816 -1131 3882 -1121
rect 4008 333 4074 389
rect 4008 -85 4074 133
rect 4008 -503 4074 -285
rect 4008 -921 4074 -703
rect 4008 -1131 4074 -1121
rect 4200 333 4266 389
rect 4200 -85 4266 133
rect 4200 -503 4266 -285
rect 4200 -921 4266 -703
rect 4200 -1131 4266 -1121
rect 4392 333 4458 389
rect 4392 -85 4458 133
rect 4392 -503 4458 -285
rect 4392 -921 4458 -703
rect 4392 -1131 4458 -1121
rect 4584 333 4650 389
rect 4584 -85 4650 133
rect 4584 -503 4650 -285
rect 4584 -921 4650 -703
rect 4584 -1131 4650 -1121
rect 4776 333 4842 389
rect 4776 -85 4842 133
rect 4776 -503 4842 -285
rect 4776 -921 4842 -703
rect 4776 -1131 4842 -1121
rect 4968 333 5034 389
rect 4968 -85 5034 133
rect 4968 -503 5034 -285
rect 4968 -921 5034 -703
rect 4968 -1131 5034 -1121
rect 5160 333 5226 389
rect 5160 -85 5226 133
rect 5160 -503 5226 -285
rect 5160 -921 5226 -703
rect 5160 -1131 5226 -1121
rect 5352 333 5418 389
rect 5352 -85 5418 133
rect 5352 -503 5418 -285
rect 5352 -921 5418 -703
rect 5352 -1131 5418 -1121
rect 5544 333 5610 389
rect 5544 -85 5610 133
rect 5544 -503 5610 -285
rect 5544 -921 5610 -703
rect 5544 -1131 5610 -1121
rect 5736 333 5802 389
rect 5736 -85 5802 133
rect 5736 -503 5802 -285
rect 5736 -921 5802 -703
rect 5736 -1131 5802 -1121
rect 5928 333 5994 389
rect 5928 -85 5994 133
rect 5928 -503 5994 -285
rect 5928 -921 5994 -703
rect 5928 -1131 5994 -1121
use sky130_fd_pr__nfet_01v8_lvt_9B2JY7  sky130_fd_pr__nfet_01v8_lvt_9B2JY7_0 ~/sky130-mpw2-fulgor/iref_ctrl_res_amp/mag
timestamp 1624020979
transform 1 0 791 0 1 -1029
box -455 -310 455 310
use sky130_fd_pr__nfet_01v8_lvt_9B2JY7  sky130_fd_pr__nfet_01v8_lvt_9B2JY7_1
timestamp 1624020979
transform 1 0 1595 0 1 -1029
box -455 -310 455 310
use sky130_fd_pr__nfet_01v8_lvt_CFLRKA  sky130_fd_pr__nfet_01v8_lvt_CFLRKA_0
timestamp 1623991863
transform 1 0 4137 0 1 956
box -2087 -519 2087 519
use sky130_fd_pr__nfet_01v8_lvt_CAF2P9  sky130_fd_pr__nfet_01v8_lvt_CAF2P9_0
timestamp 1623991863
transform 1 0 4137 0 1 -394
box -2087 -937 2087 937
<< labels >>
rlabel metal1 1164 -745 1194 -720 1 iref
rlabel metal1 356 -1340 386 -1315 1 avss1p8
rlabel metal1 2220 1481 2250 1506 1 avdd1p8
rlabel metal2 5952 522 5982 547 1 out
rlabel metal1 2020 939 2050 964 1 in
<< end >>
