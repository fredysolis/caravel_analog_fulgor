magic
tech sky130A
magscale 1 2
timestamp 1624053471
<< pwell >>
rect -16462 -24206 34360 5780
<< psubdiff >>
rect -16450 4360 -14850 4384
rect -16450 -21664 -14850 -21640
rect 32749 4360 34349 4384
rect -16450 -22594 -14851 -21664
rect 32749 -22593 34349 -21640
rect 32749 -22594 34348 -22593
rect -16450 -24194 -11039 -22594
rect 28961 -24194 34348 -22594
<< psubdiffcont >>
rect -16450 -21640 -14850 4360
rect 32749 -21640 34349 4360
rect -11039 -24194 28961 -22594
<< locali >>
rect -16450 4360 -14850 4376
rect 32749 4360 34349 4376
rect -14851 -21656 -14850 -21640
rect 34348 -21656 34349 -21640
<< viali >>
rect -16450 -21640 -14850 4360
rect 135 -119 4328 -40
rect -7307 -9814 -6904 -9752
rect -7302 -10770 -6916 -10690
rect -16450 -22594 -14851 -21640
rect 32749 -21640 34349 4360
rect 32749 -22594 34348 -21640
rect -16450 -24194 -11039 -22594
rect -11039 -24194 28961 -22594
rect 28961 -24194 34348 -22594
<< metal1 >>
rect -370 5080 -360 5680
rect 640 5614 650 5680
rect 2456 5614 2466 5680
rect 640 5182 1312 5614
rect 1560 5182 2466 5614
rect 640 5080 650 5182
rect 2456 5080 2466 5182
rect 3866 5614 3876 5680
rect 3866 5182 4100 5614
rect 3866 5080 3876 5182
rect -16456 4360 -14844 4372
rect -16456 -21634 -16450 4360
rect -16462 -24194 -16450 -21634
rect -14850 -21634 -14844 4360
rect 32743 4360 34355 4372
rect 166 166 3245 598
rect 40 -40 4361 83
rect 40 -119 135 -40
rect 4328 -119 4361 -40
rect 40 -213 4361 -119
rect 1312 -1221 2954 -213
rect 1312 -1273 2955 -1221
rect 1313 -2326 2955 -1273
rect 1313 -9453 2954 -2326
rect -6504 -9727 2954 -9453
rect -6991 -9746 2954 -9727
rect -7319 -9752 2954 -9746
rect -7319 -9814 -7307 -9752
rect -6904 -9814 2954 -9752
rect -7319 -9820 2954 -9814
rect -6991 -9828 2954 -9820
rect -6504 -9899 2954 -9828
rect -7439 -10421 -7429 -9948
rect -7166 -10421 -7156 -9948
rect -7058 -10418 -7048 -9951
rect -6795 -10418 -6785 -9951
rect -6504 -10023 -5622 -9899
rect -5632 -10420 -5622 -10023
rect -6603 -10492 -5622 -10420
rect -3065 -10023 2954 -9899
rect -3065 -10420 -3055 -10023
rect 1313 -10420 2954 -10023
rect -3065 -10492 2954 -10420
rect -8110 -10653 -7078 -10573
rect -6603 -10638 2954 -10492
rect -7010 -10684 2954 -10638
rect -7314 -10690 2954 -10684
rect -7314 -10770 -7302 -10690
rect -6916 -10770 2954 -10690
rect -7314 -10776 2954 -10770
rect -7010 -10794 2954 -10776
rect -6603 -10990 2954 -10794
rect -14850 -21640 -14839 -21634
rect -14851 -22588 -14839 -21640
rect 1313 -22588 2954 -10990
rect 32743 -22588 32749 4360
rect 34349 -21640 34355 4360
rect -14851 -22594 32749 -22588
rect 34348 -21652 34355 -21640
rect 34348 -22588 34354 -21652
rect 34348 -24194 34360 -22588
rect -16462 -24200 34360 -24194
rect 32743 -24206 34354 -24200
<< via1 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -7429 -10421 -7166 -9948
rect -7048 -10418 -6795 -9951
rect -5622 -10492 -3065 -9899
rect -16353 -24105 34174 -22697
<< metal2 >>
rect -360 5680 640 5690
rect -360 5070 640 5080
rect 2466 5680 3866 5690
rect 2466 5070 3866 5080
rect -5622 -9899 -3065 -9889
rect -7429 -9948 -7166 -9938
rect -7429 -10431 -7166 -10421
rect -7048 -9951 -6795 -9941
rect -7048 -10428 -6795 -10418
rect -5622 -10502 -3065 -10492
rect -16353 -22697 34174 -22687
rect -16353 -24115 34174 -24105
<< via2 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -7429 -10421 -7166 -9948
rect -7048 -10418 -6795 -9951
rect -5622 -10492 -3065 -9899
rect -16353 -24105 34174 -22697
<< metal3 >>
rect -370 5680 650 5685
rect -370 5080 -360 5680
rect 640 5080 650 5680
rect -370 5075 650 5080
rect 2456 5680 3876 5685
rect 2456 5080 2466 5680
rect 3866 5080 3876 5680
rect 2456 5075 3876 5080
rect -11495 -12561 -8154 -8870
rect -5655 -9894 -3064 -9027
rect -5655 -9899 -3055 -9894
rect -7439 -9948 -7156 -9943
rect -7439 -10421 -7429 -9948
rect -7166 -10421 -7156 -9948
rect -7439 -10426 -7156 -10421
rect -7058 -9951 -6785 -9946
rect -7058 -10418 -7048 -9951
rect -6795 -10418 -6785 -9951
rect -7058 -10423 -6785 -10418
rect -5655 -10492 -5622 -9899
rect -3065 -10492 -3055 -9899
rect -5655 -10497 -3055 -10492
rect -5655 -12561 -3064 -10497
rect -11495 -12710 -3064 -12561
rect -11495 -12749 -4228 -12710
rect -10301 -22692 -4228 -12749
rect 4852 -21602 9433 4898
rect 10833 -21602 14842 4898
rect 16242 -21602 20055 4898
rect 21455 -21602 25394 4898
rect 26794 -21602 31427 4898
rect 30027 -22692 31427 -21602
rect -16363 -22697 34184 -22692
rect -16363 -24105 -16353 -22697
rect 34174 -24105 34184 -22697
rect -16363 -24110 34184 -24105
<< via3 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -7429 -10421 -7166 -9948
rect -7048 -10418 -6795 -9951
<< metal4 >>
rect -10754 5680 740 5780
rect -10754 5080 -360 5680
rect 640 5080 740 5680
rect -10754 4980 740 5080
rect 2066 5680 28119 5780
rect 2066 5080 2466 5680
rect 3866 5080 28119 5680
rect 2066 4980 28119 5080
rect -7435 -9947 -7175 -7442
rect -7435 -9948 -7165 -9947
rect -7435 -10418 -7429 -9948
rect -7430 -10421 -7429 -10418
rect -7166 -10421 -7165 -9948
rect -7049 -9951 -6794 -9950
rect -7049 -10418 -7048 -9951
rect -6795 -10418 -6794 -9951
rect -7049 -10419 -6794 -10418
rect -7430 -10422 -7165 -10421
rect -7025 -11171 -6797 -10419
use sky130_fd_pr__nfet_01v8_U2JGXT  sky130_fd_pr__nfet_01v8_U2JGXT_0
timestamp 1624053471
transform 1 0 -7109 0 1 -10245
box -226 -510 226 510
use cap3_loop_filter  cap3_loop_filter_0
timestamp 1624020278
transform 1 0 -16372 0 1 -14182
box 4830 -7521 13448 3227
use res_loop_filter  res_loop_filter_2
timestamp 1624049879
transform 1 0 2956 0 1 0
box 0 0 1478 5780
use res_loop_filter  res_loop_filter_1
timestamp 1624049879
transform 1 0 1478 0 1 0
box 0 0 1478 5780
use res_loop_filter  res_loop_filter_0
timestamp 1624049879
transform 1 0 0 0 1 0
box 0 0 1478 5780
use cap1_loop_filter  cap1_loop_filter_0
timestamp 1624049879
transform 1 0 47404 0 1 20622
box -42552 -43690 -15977 -14842
use cap2_loop_filter  cap2_loop_filter_0
timestamp 1624049879
transform 1 0 -4885 0 1 288
box -8638 -9892 4299 5492
<< labels >>
rlabel pwell 1313 -22594 2954 -168 1 vss
rlabel metal4 -10754 4980 -360 5780 1 in
rlabel metal4 3866 4980 28119 5780 1 vc_pex
rlabel metal1 -8110 -10653 -7078 -10573 1 D0_cap
<< end >>
