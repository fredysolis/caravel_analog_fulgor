magic
tech sky130A
magscale 1 2
timestamp 1623991863
<< error_p >>
rect -1887 749 -1857 753
rect -1791 749 -1761 753
rect -1695 749 -1665 753
rect -1599 749 -1569 753
rect -1503 749 -1473 753
rect -1407 749 -1377 753
rect -1311 749 -1281 753
rect -1215 749 -1185 753
rect -1119 749 -1089 753
rect -1023 749 -993 753
rect -927 749 -897 753
rect -831 749 -801 753
rect -735 749 -705 753
rect -639 749 -609 753
rect -543 749 -513 753
rect -447 749 -417 753
rect -351 749 -321 753
rect -255 749 -225 753
rect -159 749 -129 753
rect -63 749 -33 753
rect 33 749 63 753
rect 129 749 159 753
rect 225 749 255 753
rect 321 749 351 753
rect 417 749 447 753
rect 513 749 543 753
rect 609 749 639 753
rect 705 749 735 753
rect 801 749 831 753
rect 897 749 927 753
rect 993 749 1023 753
rect 1089 749 1119 753
rect 1185 749 1215 753
rect 1281 749 1311 753
rect 1377 749 1407 753
rect 1473 749 1503 753
rect 1569 749 1599 753
rect 1665 749 1695 753
rect 1761 749 1791 753
rect -1887 -753 -1857 -749
rect -1791 -753 -1761 -749
rect -1695 -753 -1665 -749
rect -1599 -753 -1569 -749
rect -1503 -753 -1473 -749
rect -1407 -753 -1377 -749
rect -1311 -753 -1281 -749
rect -1215 -753 -1185 -749
rect -1119 -753 -1089 -749
rect -1023 -753 -993 -749
rect -927 -753 -897 -749
rect -831 -753 -801 -749
rect -735 -753 -705 -749
rect -639 -753 -609 -749
rect -543 -753 -513 -749
rect -447 -753 -417 -749
rect -351 -753 -321 -749
rect -255 -753 -225 -749
rect -159 -753 -129 -749
rect -63 -753 -33 -749
rect 33 -753 63 -749
rect 129 -753 159 -749
rect 225 -753 255 -749
rect 321 -753 351 -749
rect 417 -753 447 -749
rect 513 -753 543 -749
rect 609 -753 639 -749
rect 705 -753 735 -749
rect 801 -753 831 -749
rect 897 -753 927 -749
rect 993 -753 1023 -749
rect 1089 -753 1119 -749
rect 1185 -753 1215 -749
rect 1281 -753 1311 -749
rect 1377 -753 1407 -749
rect 1473 -753 1503 -749
rect 1569 -753 1599 -749
rect 1665 -753 1695 -749
rect 1761 -753 1791 -749
<< pwell >>
rect -2087 -937 2087 937
<< nmoslvt >>
rect -1887 527 -1857 727
rect -1791 527 -1761 727
rect -1695 527 -1665 727
rect -1599 527 -1569 727
rect -1503 527 -1473 727
rect -1407 527 -1377 727
rect -1311 527 -1281 727
rect -1215 527 -1185 727
rect -1119 527 -1089 727
rect -1023 527 -993 727
rect -927 527 -897 727
rect -831 527 -801 727
rect -735 527 -705 727
rect -639 527 -609 727
rect -543 527 -513 727
rect -447 527 -417 727
rect -351 527 -321 727
rect -255 527 -225 727
rect -159 527 -129 727
rect -63 527 -33 727
rect 33 527 63 727
rect 129 527 159 727
rect 225 527 255 727
rect 321 527 351 727
rect 417 527 447 727
rect 513 527 543 727
rect 609 527 639 727
rect 705 527 735 727
rect 801 527 831 727
rect 897 527 927 727
rect 993 527 1023 727
rect 1089 527 1119 727
rect 1185 527 1215 727
rect 1281 527 1311 727
rect 1377 527 1407 727
rect 1473 527 1503 727
rect 1569 527 1599 727
rect 1665 527 1695 727
rect 1761 527 1791 727
rect 1857 527 1887 727
rect -1887 109 -1857 309
rect -1791 109 -1761 309
rect -1695 109 -1665 309
rect -1599 109 -1569 309
rect -1503 109 -1473 309
rect -1407 109 -1377 309
rect -1311 109 -1281 309
rect -1215 109 -1185 309
rect -1119 109 -1089 309
rect -1023 109 -993 309
rect -927 109 -897 309
rect -831 109 -801 309
rect -735 109 -705 309
rect -639 109 -609 309
rect -543 109 -513 309
rect -447 109 -417 309
rect -351 109 -321 309
rect -255 109 -225 309
rect -159 109 -129 309
rect -63 109 -33 309
rect 33 109 63 309
rect 129 109 159 309
rect 225 109 255 309
rect 321 109 351 309
rect 417 109 447 309
rect 513 109 543 309
rect 609 109 639 309
rect 705 109 735 309
rect 801 109 831 309
rect 897 109 927 309
rect 993 109 1023 309
rect 1089 109 1119 309
rect 1185 109 1215 309
rect 1281 109 1311 309
rect 1377 109 1407 309
rect 1473 109 1503 309
rect 1569 109 1599 309
rect 1665 109 1695 309
rect 1761 109 1791 309
rect 1857 109 1887 309
rect -1887 -309 -1857 -109
rect -1791 -309 -1761 -109
rect -1695 -309 -1665 -109
rect -1599 -309 -1569 -109
rect -1503 -309 -1473 -109
rect -1407 -309 -1377 -109
rect -1311 -309 -1281 -109
rect -1215 -309 -1185 -109
rect -1119 -309 -1089 -109
rect -1023 -309 -993 -109
rect -927 -309 -897 -109
rect -831 -309 -801 -109
rect -735 -309 -705 -109
rect -639 -309 -609 -109
rect -543 -309 -513 -109
rect -447 -309 -417 -109
rect -351 -309 -321 -109
rect -255 -309 -225 -109
rect -159 -309 -129 -109
rect -63 -309 -33 -109
rect 33 -309 63 -109
rect 129 -309 159 -109
rect 225 -309 255 -109
rect 321 -309 351 -109
rect 417 -309 447 -109
rect 513 -309 543 -109
rect 609 -309 639 -109
rect 705 -309 735 -109
rect 801 -309 831 -109
rect 897 -309 927 -109
rect 993 -309 1023 -109
rect 1089 -309 1119 -109
rect 1185 -309 1215 -109
rect 1281 -309 1311 -109
rect 1377 -309 1407 -109
rect 1473 -309 1503 -109
rect 1569 -309 1599 -109
rect 1665 -309 1695 -109
rect 1761 -309 1791 -109
rect 1857 -309 1887 -109
rect -1887 -727 -1857 -527
rect -1791 -727 -1761 -527
rect -1695 -727 -1665 -527
rect -1599 -727 -1569 -527
rect -1503 -727 -1473 -527
rect -1407 -727 -1377 -527
rect -1311 -727 -1281 -527
rect -1215 -727 -1185 -527
rect -1119 -727 -1089 -527
rect -1023 -727 -993 -527
rect -927 -727 -897 -527
rect -831 -727 -801 -527
rect -735 -727 -705 -527
rect -639 -727 -609 -527
rect -543 -727 -513 -527
rect -447 -727 -417 -527
rect -351 -727 -321 -527
rect -255 -727 -225 -527
rect -159 -727 -129 -527
rect -63 -727 -33 -527
rect 33 -727 63 -527
rect 129 -727 159 -527
rect 225 -727 255 -527
rect 321 -727 351 -527
rect 417 -727 447 -527
rect 513 -727 543 -527
rect 609 -727 639 -527
rect 705 -727 735 -527
rect 801 -727 831 -527
rect 897 -727 927 -527
rect 993 -727 1023 -527
rect 1089 -727 1119 -527
rect 1185 -727 1215 -527
rect 1281 -727 1311 -527
rect 1377 -727 1407 -527
rect 1473 -727 1503 -527
rect 1569 -727 1599 -527
rect 1665 -727 1695 -527
rect 1761 -727 1791 -527
rect 1857 -727 1887 -527
<< ndiff >>
rect -1949 715 -1887 727
rect -1949 539 -1937 715
rect -1903 539 -1887 715
rect -1949 527 -1887 539
rect -1857 715 -1791 727
rect -1857 539 -1841 715
rect -1807 539 -1791 715
rect -1857 527 -1791 539
rect -1761 715 -1695 727
rect -1761 539 -1745 715
rect -1711 539 -1695 715
rect -1761 527 -1695 539
rect -1665 715 -1599 727
rect -1665 539 -1649 715
rect -1615 539 -1599 715
rect -1665 527 -1599 539
rect -1569 715 -1503 727
rect -1569 539 -1553 715
rect -1519 539 -1503 715
rect -1569 527 -1503 539
rect -1473 715 -1407 727
rect -1473 539 -1457 715
rect -1423 539 -1407 715
rect -1473 527 -1407 539
rect -1377 715 -1311 727
rect -1377 539 -1361 715
rect -1327 539 -1311 715
rect -1377 527 -1311 539
rect -1281 715 -1215 727
rect -1281 539 -1265 715
rect -1231 539 -1215 715
rect -1281 527 -1215 539
rect -1185 715 -1119 727
rect -1185 539 -1169 715
rect -1135 539 -1119 715
rect -1185 527 -1119 539
rect -1089 715 -1023 727
rect -1089 539 -1073 715
rect -1039 539 -1023 715
rect -1089 527 -1023 539
rect -993 715 -927 727
rect -993 539 -977 715
rect -943 539 -927 715
rect -993 527 -927 539
rect -897 715 -831 727
rect -897 539 -881 715
rect -847 539 -831 715
rect -897 527 -831 539
rect -801 715 -735 727
rect -801 539 -785 715
rect -751 539 -735 715
rect -801 527 -735 539
rect -705 715 -639 727
rect -705 539 -689 715
rect -655 539 -639 715
rect -705 527 -639 539
rect -609 715 -543 727
rect -609 539 -593 715
rect -559 539 -543 715
rect -609 527 -543 539
rect -513 715 -447 727
rect -513 539 -497 715
rect -463 539 -447 715
rect -513 527 -447 539
rect -417 715 -351 727
rect -417 539 -401 715
rect -367 539 -351 715
rect -417 527 -351 539
rect -321 715 -255 727
rect -321 539 -305 715
rect -271 539 -255 715
rect -321 527 -255 539
rect -225 715 -159 727
rect -225 539 -209 715
rect -175 539 -159 715
rect -225 527 -159 539
rect -129 715 -63 727
rect -129 539 -113 715
rect -79 539 -63 715
rect -129 527 -63 539
rect -33 715 33 727
rect -33 539 -17 715
rect 17 539 33 715
rect -33 527 33 539
rect 63 715 129 727
rect 63 539 79 715
rect 113 539 129 715
rect 63 527 129 539
rect 159 715 225 727
rect 159 539 175 715
rect 209 539 225 715
rect 159 527 225 539
rect 255 715 321 727
rect 255 539 271 715
rect 305 539 321 715
rect 255 527 321 539
rect 351 715 417 727
rect 351 539 367 715
rect 401 539 417 715
rect 351 527 417 539
rect 447 715 513 727
rect 447 539 463 715
rect 497 539 513 715
rect 447 527 513 539
rect 543 715 609 727
rect 543 539 559 715
rect 593 539 609 715
rect 543 527 609 539
rect 639 715 705 727
rect 639 539 655 715
rect 689 539 705 715
rect 639 527 705 539
rect 735 715 801 727
rect 735 539 751 715
rect 785 539 801 715
rect 735 527 801 539
rect 831 715 897 727
rect 831 539 847 715
rect 881 539 897 715
rect 831 527 897 539
rect 927 715 993 727
rect 927 539 943 715
rect 977 539 993 715
rect 927 527 993 539
rect 1023 715 1089 727
rect 1023 539 1039 715
rect 1073 539 1089 715
rect 1023 527 1089 539
rect 1119 715 1185 727
rect 1119 539 1135 715
rect 1169 539 1185 715
rect 1119 527 1185 539
rect 1215 715 1281 727
rect 1215 539 1231 715
rect 1265 539 1281 715
rect 1215 527 1281 539
rect 1311 715 1377 727
rect 1311 539 1327 715
rect 1361 539 1377 715
rect 1311 527 1377 539
rect 1407 715 1473 727
rect 1407 539 1423 715
rect 1457 539 1473 715
rect 1407 527 1473 539
rect 1503 715 1569 727
rect 1503 539 1519 715
rect 1553 539 1569 715
rect 1503 527 1569 539
rect 1599 715 1665 727
rect 1599 539 1615 715
rect 1649 539 1665 715
rect 1599 527 1665 539
rect 1695 715 1761 727
rect 1695 539 1711 715
rect 1745 539 1761 715
rect 1695 527 1761 539
rect 1791 715 1857 727
rect 1791 539 1807 715
rect 1841 539 1857 715
rect 1791 527 1857 539
rect 1887 715 1949 727
rect 1887 539 1903 715
rect 1937 539 1949 715
rect 1887 527 1949 539
rect -1949 297 -1887 309
rect -1949 121 -1937 297
rect -1903 121 -1887 297
rect -1949 109 -1887 121
rect -1857 297 -1791 309
rect -1857 121 -1841 297
rect -1807 121 -1791 297
rect -1857 109 -1791 121
rect -1761 297 -1695 309
rect -1761 121 -1745 297
rect -1711 121 -1695 297
rect -1761 109 -1695 121
rect -1665 297 -1599 309
rect -1665 121 -1649 297
rect -1615 121 -1599 297
rect -1665 109 -1599 121
rect -1569 297 -1503 309
rect -1569 121 -1553 297
rect -1519 121 -1503 297
rect -1569 109 -1503 121
rect -1473 297 -1407 309
rect -1473 121 -1457 297
rect -1423 121 -1407 297
rect -1473 109 -1407 121
rect -1377 297 -1311 309
rect -1377 121 -1361 297
rect -1327 121 -1311 297
rect -1377 109 -1311 121
rect -1281 297 -1215 309
rect -1281 121 -1265 297
rect -1231 121 -1215 297
rect -1281 109 -1215 121
rect -1185 297 -1119 309
rect -1185 121 -1169 297
rect -1135 121 -1119 297
rect -1185 109 -1119 121
rect -1089 297 -1023 309
rect -1089 121 -1073 297
rect -1039 121 -1023 297
rect -1089 109 -1023 121
rect -993 297 -927 309
rect -993 121 -977 297
rect -943 121 -927 297
rect -993 109 -927 121
rect -897 297 -831 309
rect -897 121 -881 297
rect -847 121 -831 297
rect -897 109 -831 121
rect -801 297 -735 309
rect -801 121 -785 297
rect -751 121 -735 297
rect -801 109 -735 121
rect -705 297 -639 309
rect -705 121 -689 297
rect -655 121 -639 297
rect -705 109 -639 121
rect -609 297 -543 309
rect -609 121 -593 297
rect -559 121 -543 297
rect -609 109 -543 121
rect -513 297 -447 309
rect -513 121 -497 297
rect -463 121 -447 297
rect -513 109 -447 121
rect -417 297 -351 309
rect -417 121 -401 297
rect -367 121 -351 297
rect -417 109 -351 121
rect -321 297 -255 309
rect -321 121 -305 297
rect -271 121 -255 297
rect -321 109 -255 121
rect -225 297 -159 309
rect -225 121 -209 297
rect -175 121 -159 297
rect -225 109 -159 121
rect -129 297 -63 309
rect -129 121 -113 297
rect -79 121 -63 297
rect -129 109 -63 121
rect -33 297 33 309
rect -33 121 -17 297
rect 17 121 33 297
rect -33 109 33 121
rect 63 297 129 309
rect 63 121 79 297
rect 113 121 129 297
rect 63 109 129 121
rect 159 297 225 309
rect 159 121 175 297
rect 209 121 225 297
rect 159 109 225 121
rect 255 297 321 309
rect 255 121 271 297
rect 305 121 321 297
rect 255 109 321 121
rect 351 297 417 309
rect 351 121 367 297
rect 401 121 417 297
rect 351 109 417 121
rect 447 297 513 309
rect 447 121 463 297
rect 497 121 513 297
rect 447 109 513 121
rect 543 297 609 309
rect 543 121 559 297
rect 593 121 609 297
rect 543 109 609 121
rect 639 297 705 309
rect 639 121 655 297
rect 689 121 705 297
rect 639 109 705 121
rect 735 297 801 309
rect 735 121 751 297
rect 785 121 801 297
rect 735 109 801 121
rect 831 297 897 309
rect 831 121 847 297
rect 881 121 897 297
rect 831 109 897 121
rect 927 297 993 309
rect 927 121 943 297
rect 977 121 993 297
rect 927 109 993 121
rect 1023 297 1089 309
rect 1023 121 1039 297
rect 1073 121 1089 297
rect 1023 109 1089 121
rect 1119 297 1185 309
rect 1119 121 1135 297
rect 1169 121 1185 297
rect 1119 109 1185 121
rect 1215 297 1281 309
rect 1215 121 1231 297
rect 1265 121 1281 297
rect 1215 109 1281 121
rect 1311 297 1377 309
rect 1311 121 1327 297
rect 1361 121 1377 297
rect 1311 109 1377 121
rect 1407 297 1473 309
rect 1407 121 1423 297
rect 1457 121 1473 297
rect 1407 109 1473 121
rect 1503 297 1569 309
rect 1503 121 1519 297
rect 1553 121 1569 297
rect 1503 109 1569 121
rect 1599 297 1665 309
rect 1599 121 1615 297
rect 1649 121 1665 297
rect 1599 109 1665 121
rect 1695 297 1761 309
rect 1695 121 1711 297
rect 1745 121 1761 297
rect 1695 109 1761 121
rect 1791 297 1857 309
rect 1791 121 1807 297
rect 1841 121 1857 297
rect 1791 109 1857 121
rect 1887 297 1949 309
rect 1887 121 1903 297
rect 1937 121 1949 297
rect 1887 109 1949 121
rect -1949 -121 -1887 -109
rect -1949 -297 -1937 -121
rect -1903 -297 -1887 -121
rect -1949 -309 -1887 -297
rect -1857 -121 -1791 -109
rect -1857 -297 -1841 -121
rect -1807 -297 -1791 -121
rect -1857 -309 -1791 -297
rect -1761 -121 -1695 -109
rect -1761 -297 -1745 -121
rect -1711 -297 -1695 -121
rect -1761 -309 -1695 -297
rect -1665 -121 -1599 -109
rect -1665 -297 -1649 -121
rect -1615 -297 -1599 -121
rect -1665 -309 -1599 -297
rect -1569 -121 -1503 -109
rect -1569 -297 -1553 -121
rect -1519 -297 -1503 -121
rect -1569 -309 -1503 -297
rect -1473 -121 -1407 -109
rect -1473 -297 -1457 -121
rect -1423 -297 -1407 -121
rect -1473 -309 -1407 -297
rect -1377 -121 -1311 -109
rect -1377 -297 -1361 -121
rect -1327 -297 -1311 -121
rect -1377 -309 -1311 -297
rect -1281 -121 -1215 -109
rect -1281 -297 -1265 -121
rect -1231 -297 -1215 -121
rect -1281 -309 -1215 -297
rect -1185 -121 -1119 -109
rect -1185 -297 -1169 -121
rect -1135 -297 -1119 -121
rect -1185 -309 -1119 -297
rect -1089 -121 -1023 -109
rect -1089 -297 -1073 -121
rect -1039 -297 -1023 -121
rect -1089 -309 -1023 -297
rect -993 -121 -927 -109
rect -993 -297 -977 -121
rect -943 -297 -927 -121
rect -993 -309 -927 -297
rect -897 -121 -831 -109
rect -897 -297 -881 -121
rect -847 -297 -831 -121
rect -897 -309 -831 -297
rect -801 -121 -735 -109
rect -801 -297 -785 -121
rect -751 -297 -735 -121
rect -801 -309 -735 -297
rect -705 -121 -639 -109
rect -705 -297 -689 -121
rect -655 -297 -639 -121
rect -705 -309 -639 -297
rect -609 -121 -543 -109
rect -609 -297 -593 -121
rect -559 -297 -543 -121
rect -609 -309 -543 -297
rect -513 -121 -447 -109
rect -513 -297 -497 -121
rect -463 -297 -447 -121
rect -513 -309 -447 -297
rect -417 -121 -351 -109
rect -417 -297 -401 -121
rect -367 -297 -351 -121
rect -417 -309 -351 -297
rect -321 -121 -255 -109
rect -321 -297 -305 -121
rect -271 -297 -255 -121
rect -321 -309 -255 -297
rect -225 -121 -159 -109
rect -225 -297 -209 -121
rect -175 -297 -159 -121
rect -225 -309 -159 -297
rect -129 -121 -63 -109
rect -129 -297 -113 -121
rect -79 -297 -63 -121
rect -129 -309 -63 -297
rect -33 -121 33 -109
rect -33 -297 -17 -121
rect 17 -297 33 -121
rect -33 -309 33 -297
rect 63 -121 129 -109
rect 63 -297 79 -121
rect 113 -297 129 -121
rect 63 -309 129 -297
rect 159 -121 225 -109
rect 159 -297 175 -121
rect 209 -297 225 -121
rect 159 -309 225 -297
rect 255 -121 321 -109
rect 255 -297 271 -121
rect 305 -297 321 -121
rect 255 -309 321 -297
rect 351 -121 417 -109
rect 351 -297 367 -121
rect 401 -297 417 -121
rect 351 -309 417 -297
rect 447 -121 513 -109
rect 447 -297 463 -121
rect 497 -297 513 -121
rect 447 -309 513 -297
rect 543 -121 609 -109
rect 543 -297 559 -121
rect 593 -297 609 -121
rect 543 -309 609 -297
rect 639 -121 705 -109
rect 639 -297 655 -121
rect 689 -297 705 -121
rect 639 -309 705 -297
rect 735 -121 801 -109
rect 735 -297 751 -121
rect 785 -297 801 -121
rect 735 -309 801 -297
rect 831 -121 897 -109
rect 831 -297 847 -121
rect 881 -297 897 -121
rect 831 -309 897 -297
rect 927 -121 993 -109
rect 927 -297 943 -121
rect 977 -297 993 -121
rect 927 -309 993 -297
rect 1023 -121 1089 -109
rect 1023 -297 1039 -121
rect 1073 -297 1089 -121
rect 1023 -309 1089 -297
rect 1119 -121 1185 -109
rect 1119 -297 1135 -121
rect 1169 -297 1185 -121
rect 1119 -309 1185 -297
rect 1215 -121 1281 -109
rect 1215 -297 1231 -121
rect 1265 -297 1281 -121
rect 1215 -309 1281 -297
rect 1311 -121 1377 -109
rect 1311 -297 1327 -121
rect 1361 -297 1377 -121
rect 1311 -309 1377 -297
rect 1407 -121 1473 -109
rect 1407 -297 1423 -121
rect 1457 -297 1473 -121
rect 1407 -309 1473 -297
rect 1503 -121 1569 -109
rect 1503 -297 1519 -121
rect 1553 -297 1569 -121
rect 1503 -309 1569 -297
rect 1599 -121 1665 -109
rect 1599 -297 1615 -121
rect 1649 -297 1665 -121
rect 1599 -309 1665 -297
rect 1695 -121 1761 -109
rect 1695 -297 1711 -121
rect 1745 -297 1761 -121
rect 1695 -309 1761 -297
rect 1791 -121 1857 -109
rect 1791 -297 1807 -121
rect 1841 -297 1857 -121
rect 1791 -309 1857 -297
rect 1887 -121 1949 -109
rect 1887 -297 1903 -121
rect 1937 -297 1949 -121
rect 1887 -309 1949 -297
rect -1949 -539 -1887 -527
rect -1949 -715 -1937 -539
rect -1903 -715 -1887 -539
rect -1949 -727 -1887 -715
rect -1857 -539 -1791 -527
rect -1857 -715 -1841 -539
rect -1807 -715 -1791 -539
rect -1857 -727 -1791 -715
rect -1761 -539 -1695 -527
rect -1761 -715 -1745 -539
rect -1711 -715 -1695 -539
rect -1761 -727 -1695 -715
rect -1665 -539 -1599 -527
rect -1665 -715 -1649 -539
rect -1615 -715 -1599 -539
rect -1665 -727 -1599 -715
rect -1569 -539 -1503 -527
rect -1569 -715 -1553 -539
rect -1519 -715 -1503 -539
rect -1569 -727 -1503 -715
rect -1473 -539 -1407 -527
rect -1473 -715 -1457 -539
rect -1423 -715 -1407 -539
rect -1473 -727 -1407 -715
rect -1377 -539 -1311 -527
rect -1377 -715 -1361 -539
rect -1327 -715 -1311 -539
rect -1377 -727 -1311 -715
rect -1281 -539 -1215 -527
rect -1281 -715 -1265 -539
rect -1231 -715 -1215 -539
rect -1281 -727 -1215 -715
rect -1185 -539 -1119 -527
rect -1185 -715 -1169 -539
rect -1135 -715 -1119 -539
rect -1185 -727 -1119 -715
rect -1089 -539 -1023 -527
rect -1089 -715 -1073 -539
rect -1039 -715 -1023 -539
rect -1089 -727 -1023 -715
rect -993 -539 -927 -527
rect -993 -715 -977 -539
rect -943 -715 -927 -539
rect -993 -727 -927 -715
rect -897 -539 -831 -527
rect -897 -715 -881 -539
rect -847 -715 -831 -539
rect -897 -727 -831 -715
rect -801 -539 -735 -527
rect -801 -715 -785 -539
rect -751 -715 -735 -539
rect -801 -727 -735 -715
rect -705 -539 -639 -527
rect -705 -715 -689 -539
rect -655 -715 -639 -539
rect -705 -727 -639 -715
rect -609 -539 -543 -527
rect -609 -715 -593 -539
rect -559 -715 -543 -539
rect -609 -727 -543 -715
rect -513 -539 -447 -527
rect -513 -715 -497 -539
rect -463 -715 -447 -539
rect -513 -727 -447 -715
rect -417 -539 -351 -527
rect -417 -715 -401 -539
rect -367 -715 -351 -539
rect -417 -727 -351 -715
rect -321 -539 -255 -527
rect -321 -715 -305 -539
rect -271 -715 -255 -539
rect -321 -727 -255 -715
rect -225 -539 -159 -527
rect -225 -715 -209 -539
rect -175 -715 -159 -539
rect -225 -727 -159 -715
rect -129 -539 -63 -527
rect -129 -715 -113 -539
rect -79 -715 -63 -539
rect -129 -727 -63 -715
rect -33 -539 33 -527
rect -33 -715 -17 -539
rect 17 -715 33 -539
rect -33 -727 33 -715
rect 63 -539 129 -527
rect 63 -715 79 -539
rect 113 -715 129 -539
rect 63 -727 129 -715
rect 159 -539 225 -527
rect 159 -715 175 -539
rect 209 -715 225 -539
rect 159 -727 225 -715
rect 255 -539 321 -527
rect 255 -715 271 -539
rect 305 -715 321 -539
rect 255 -727 321 -715
rect 351 -539 417 -527
rect 351 -715 367 -539
rect 401 -715 417 -539
rect 351 -727 417 -715
rect 447 -539 513 -527
rect 447 -715 463 -539
rect 497 -715 513 -539
rect 447 -727 513 -715
rect 543 -539 609 -527
rect 543 -715 559 -539
rect 593 -715 609 -539
rect 543 -727 609 -715
rect 639 -539 705 -527
rect 639 -715 655 -539
rect 689 -715 705 -539
rect 639 -727 705 -715
rect 735 -539 801 -527
rect 735 -715 751 -539
rect 785 -715 801 -539
rect 735 -727 801 -715
rect 831 -539 897 -527
rect 831 -715 847 -539
rect 881 -715 897 -539
rect 831 -727 897 -715
rect 927 -539 993 -527
rect 927 -715 943 -539
rect 977 -715 993 -539
rect 927 -727 993 -715
rect 1023 -539 1089 -527
rect 1023 -715 1039 -539
rect 1073 -715 1089 -539
rect 1023 -727 1089 -715
rect 1119 -539 1185 -527
rect 1119 -715 1135 -539
rect 1169 -715 1185 -539
rect 1119 -727 1185 -715
rect 1215 -539 1281 -527
rect 1215 -715 1231 -539
rect 1265 -715 1281 -539
rect 1215 -727 1281 -715
rect 1311 -539 1377 -527
rect 1311 -715 1327 -539
rect 1361 -715 1377 -539
rect 1311 -727 1377 -715
rect 1407 -539 1473 -527
rect 1407 -715 1423 -539
rect 1457 -715 1473 -539
rect 1407 -727 1473 -715
rect 1503 -539 1569 -527
rect 1503 -715 1519 -539
rect 1553 -715 1569 -539
rect 1503 -727 1569 -715
rect 1599 -539 1665 -527
rect 1599 -715 1615 -539
rect 1649 -715 1665 -539
rect 1599 -727 1665 -715
rect 1695 -539 1761 -527
rect 1695 -715 1711 -539
rect 1745 -715 1761 -539
rect 1695 -727 1761 -715
rect 1791 -539 1857 -527
rect 1791 -715 1807 -539
rect 1841 -715 1857 -539
rect 1791 -727 1857 -715
rect 1887 -539 1949 -527
rect 1887 -715 1903 -539
rect 1937 -715 1949 -539
rect 1887 -727 1949 -715
<< ndiffc >>
rect -1937 539 -1903 715
rect -1841 539 -1807 715
rect -1745 539 -1711 715
rect -1649 539 -1615 715
rect -1553 539 -1519 715
rect -1457 539 -1423 715
rect -1361 539 -1327 715
rect -1265 539 -1231 715
rect -1169 539 -1135 715
rect -1073 539 -1039 715
rect -977 539 -943 715
rect -881 539 -847 715
rect -785 539 -751 715
rect -689 539 -655 715
rect -593 539 -559 715
rect -497 539 -463 715
rect -401 539 -367 715
rect -305 539 -271 715
rect -209 539 -175 715
rect -113 539 -79 715
rect -17 539 17 715
rect 79 539 113 715
rect 175 539 209 715
rect 271 539 305 715
rect 367 539 401 715
rect 463 539 497 715
rect 559 539 593 715
rect 655 539 689 715
rect 751 539 785 715
rect 847 539 881 715
rect 943 539 977 715
rect 1039 539 1073 715
rect 1135 539 1169 715
rect 1231 539 1265 715
rect 1327 539 1361 715
rect 1423 539 1457 715
rect 1519 539 1553 715
rect 1615 539 1649 715
rect 1711 539 1745 715
rect 1807 539 1841 715
rect 1903 539 1937 715
rect -1937 121 -1903 297
rect -1841 121 -1807 297
rect -1745 121 -1711 297
rect -1649 121 -1615 297
rect -1553 121 -1519 297
rect -1457 121 -1423 297
rect -1361 121 -1327 297
rect -1265 121 -1231 297
rect -1169 121 -1135 297
rect -1073 121 -1039 297
rect -977 121 -943 297
rect -881 121 -847 297
rect -785 121 -751 297
rect -689 121 -655 297
rect -593 121 -559 297
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect 559 121 593 297
rect 655 121 689 297
rect 751 121 785 297
rect 847 121 881 297
rect 943 121 977 297
rect 1039 121 1073 297
rect 1135 121 1169 297
rect 1231 121 1265 297
rect 1327 121 1361 297
rect 1423 121 1457 297
rect 1519 121 1553 297
rect 1615 121 1649 297
rect 1711 121 1745 297
rect 1807 121 1841 297
rect 1903 121 1937 297
rect -1937 -297 -1903 -121
rect -1841 -297 -1807 -121
rect -1745 -297 -1711 -121
rect -1649 -297 -1615 -121
rect -1553 -297 -1519 -121
rect -1457 -297 -1423 -121
rect -1361 -297 -1327 -121
rect -1265 -297 -1231 -121
rect -1169 -297 -1135 -121
rect -1073 -297 -1039 -121
rect -977 -297 -943 -121
rect -881 -297 -847 -121
rect -785 -297 -751 -121
rect -689 -297 -655 -121
rect -593 -297 -559 -121
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect 559 -297 593 -121
rect 655 -297 689 -121
rect 751 -297 785 -121
rect 847 -297 881 -121
rect 943 -297 977 -121
rect 1039 -297 1073 -121
rect 1135 -297 1169 -121
rect 1231 -297 1265 -121
rect 1327 -297 1361 -121
rect 1423 -297 1457 -121
rect 1519 -297 1553 -121
rect 1615 -297 1649 -121
rect 1711 -297 1745 -121
rect 1807 -297 1841 -121
rect 1903 -297 1937 -121
rect -1937 -715 -1903 -539
rect -1841 -715 -1807 -539
rect -1745 -715 -1711 -539
rect -1649 -715 -1615 -539
rect -1553 -715 -1519 -539
rect -1457 -715 -1423 -539
rect -1361 -715 -1327 -539
rect -1265 -715 -1231 -539
rect -1169 -715 -1135 -539
rect -1073 -715 -1039 -539
rect -977 -715 -943 -539
rect -881 -715 -847 -539
rect -785 -715 -751 -539
rect -689 -715 -655 -539
rect -593 -715 -559 -539
rect -497 -715 -463 -539
rect -401 -715 -367 -539
rect -305 -715 -271 -539
rect -209 -715 -175 -539
rect -113 -715 -79 -539
rect -17 -715 17 -539
rect 79 -715 113 -539
rect 175 -715 209 -539
rect 271 -715 305 -539
rect 367 -715 401 -539
rect 463 -715 497 -539
rect 559 -715 593 -539
rect 655 -715 689 -539
rect 751 -715 785 -539
rect 847 -715 881 -539
rect 943 -715 977 -539
rect 1039 -715 1073 -539
rect 1135 -715 1169 -539
rect 1231 -715 1265 -539
rect 1327 -715 1361 -539
rect 1423 -715 1457 -539
rect 1519 -715 1553 -539
rect 1615 -715 1649 -539
rect 1711 -715 1745 -539
rect 1807 -715 1841 -539
rect 1903 -715 1937 -539
<< psubdiff >>
rect -2051 867 -1955 901
rect 1955 867 2051 901
rect 2017 805 2051 867
rect 2017 -867 2051 -805
rect -2051 -901 -1955 -867
rect 1955 -901 2051 -867
<< psubdiffcont >>
rect -1955 867 1955 901
rect 2017 -805 2051 805
rect -1955 -901 1955 -867
<< poly >>
rect -1887 727 -1857 749
rect -1791 727 -1761 749
rect -1695 727 -1665 749
rect -1599 727 -1569 749
rect -1503 727 -1473 749
rect -1407 727 -1377 749
rect -1311 727 -1281 749
rect -1215 727 -1185 749
rect -1119 727 -1089 749
rect -1023 727 -993 749
rect -927 727 -897 749
rect -831 727 -801 749
rect -735 727 -705 749
rect -639 727 -609 749
rect -543 727 -513 749
rect -447 727 -417 749
rect -351 727 -321 749
rect -255 727 -225 749
rect -159 727 -129 749
rect -63 727 -33 749
rect 33 727 63 749
rect 129 727 159 749
rect 225 727 255 749
rect 321 727 351 749
rect 417 727 447 749
rect 513 727 543 749
rect 609 727 639 749
rect 705 727 735 749
rect 801 727 831 749
rect 897 727 927 749
rect 993 727 1023 749
rect 1089 727 1119 749
rect 1185 727 1215 749
rect 1281 727 1311 749
rect 1377 727 1407 749
rect 1473 727 1503 749
rect 1569 727 1599 749
rect 1665 727 1695 749
rect 1761 727 1791 749
rect 1857 727 1887 753
rect -1887 505 -1857 527
rect -1791 505 -1761 527
rect -1695 505 -1665 527
rect -1599 505 -1569 527
rect -1503 505 -1473 527
rect -1407 505 -1377 527
rect -1311 505 -1281 527
rect -1215 505 -1185 527
rect -1119 505 -1089 527
rect -1023 505 -993 527
rect -927 505 -897 527
rect -831 505 -801 527
rect -735 505 -705 527
rect -639 505 -609 527
rect -543 505 -513 527
rect -447 505 -417 527
rect -351 505 -321 527
rect -255 505 -225 527
rect -159 505 -129 527
rect -63 505 -33 527
rect 33 505 63 527
rect 129 505 159 527
rect 225 505 255 527
rect 321 505 351 527
rect 417 505 447 527
rect 513 505 543 527
rect 609 505 639 527
rect 705 505 735 527
rect 801 505 831 527
rect 897 505 927 527
rect 993 505 1023 527
rect 1089 505 1119 527
rect 1185 505 1215 527
rect 1281 505 1311 527
rect 1377 505 1407 527
rect 1473 505 1503 527
rect 1569 505 1599 527
rect 1665 505 1695 527
rect 1761 505 1791 527
rect 1857 505 1887 527
rect -1904 331 1906 505
rect -1887 309 -1857 331
rect -1791 309 -1761 331
rect -1695 309 -1665 331
rect -1599 309 -1569 331
rect -1503 309 -1473 331
rect -1407 309 -1377 331
rect -1311 309 -1281 331
rect -1215 309 -1185 331
rect -1119 309 -1089 331
rect -1023 309 -993 331
rect -927 309 -897 331
rect -831 309 -801 331
rect -735 309 -705 331
rect -639 309 -609 331
rect -543 309 -513 331
rect -447 309 -417 331
rect -351 309 -321 331
rect -255 309 -225 331
rect -159 309 -129 331
rect -63 309 -33 331
rect 33 309 63 331
rect 129 309 159 331
rect 225 309 255 331
rect 321 309 351 331
rect 417 309 447 331
rect 513 309 543 331
rect 609 309 639 331
rect 705 309 735 331
rect 801 309 831 331
rect 897 309 927 331
rect 993 309 1023 331
rect 1089 309 1119 331
rect 1185 309 1215 331
rect 1281 309 1311 331
rect 1377 309 1407 331
rect 1473 309 1503 331
rect 1569 309 1599 331
rect 1665 309 1695 331
rect 1761 309 1791 331
rect 1857 309 1887 331
rect -1887 87 -1857 109
rect -1791 87 -1761 109
rect -1695 87 -1665 109
rect -1599 87 -1569 109
rect -1503 87 -1473 109
rect -1407 87 -1377 109
rect -1311 87 -1281 109
rect -1215 87 -1185 109
rect -1119 87 -1089 109
rect -1023 87 -993 109
rect -927 87 -897 109
rect -831 87 -801 109
rect -735 87 -705 109
rect -639 87 -609 109
rect -543 87 -513 109
rect -447 87 -417 109
rect -351 87 -321 109
rect -255 87 -225 109
rect -159 87 -129 109
rect -63 87 -33 109
rect 33 87 63 109
rect 129 87 159 109
rect 225 87 255 109
rect 321 87 351 109
rect 417 87 447 109
rect 513 87 543 109
rect 609 87 639 109
rect 705 87 735 109
rect 801 87 831 109
rect 897 87 927 109
rect 993 87 1023 109
rect 1089 87 1119 109
rect 1185 87 1215 109
rect 1281 87 1311 109
rect 1377 87 1407 109
rect 1473 87 1503 109
rect 1569 87 1599 109
rect 1665 87 1695 109
rect 1761 87 1791 109
rect 1857 87 1887 109
rect -1905 -87 1905 87
rect -1887 -109 -1857 -87
rect -1791 -109 -1761 -87
rect -1695 -109 -1665 -87
rect -1599 -109 -1569 -87
rect -1503 -109 -1473 -87
rect -1407 -109 -1377 -87
rect -1311 -109 -1281 -87
rect -1215 -109 -1185 -87
rect -1119 -109 -1089 -87
rect -1023 -109 -993 -87
rect -927 -109 -897 -87
rect -831 -109 -801 -87
rect -735 -109 -705 -87
rect -639 -109 -609 -87
rect -543 -109 -513 -87
rect -447 -109 -417 -87
rect -351 -109 -321 -87
rect -255 -109 -225 -87
rect -159 -109 -129 -87
rect -63 -109 -33 -87
rect 33 -109 63 -87
rect 129 -109 159 -87
rect 225 -109 255 -87
rect 321 -109 351 -87
rect 417 -109 447 -87
rect 513 -109 543 -87
rect 609 -109 639 -87
rect 705 -109 735 -87
rect 801 -109 831 -87
rect 897 -109 927 -87
rect 993 -109 1023 -87
rect 1089 -109 1119 -87
rect 1185 -109 1215 -87
rect 1281 -109 1311 -87
rect 1377 -109 1407 -87
rect 1473 -109 1503 -87
rect 1569 -109 1599 -87
rect 1665 -109 1695 -87
rect 1761 -109 1791 -87
rect 1857 -109 1887 -87
rect -1887 -331 -1857 -309
rect -1791 -331 -1761 -309
rect -1695 -331 -1665 -309
rect -1599 -331 -1569 -309
rect -1503 -331 -1473 -309
rect -1407 -331 -1377 -309
rect -1311 -331 -1281 -309
rect -1215 -331 -1185 -309
rect -1119 -331 -1089 -309
rect -1023 -331 -993 -309
rect -927 -331 -897 -309
rect -831 -331 -801 -309
rect -735 -331 -705 -309
rect -639 -331 -609 -309
rect -543 -331 -513 -309
rect -447 -331 -417 -309
rect -351 -331 -321 -309
rect -255 -331 -225 -309
rect -159 -331 -129 -309
rect -63 -331 -33 -309
rect 33 -331 63 -309
rect 129 -331 159 -309
rect 225 -331 255 -309
rect 321 -331 351 -309
rect 417 -331 447 -309
rect 513 -331 543 -309
rect 609 -331 639 -309
rect 705 -331 735 -309
rect 801 -331 831 -309
rect 897 -331 927 -309
rect 993 -331 1023 -309
rect 1089 -331 1119 -309
rect 1185 -331 1215 -309
rect 1281 -331 1311 -309
rect 1377 -331 1407 -309
rect 1473 -331 1503 -309
rect 1569 -331 1599 -309
rect 1665 -331 1695 -309
rect 1761 -331 1791 -309
rect 1857 -331 1887 -309
rect -1905 -505 1905 -331
rect -1887 -527 -1857 -505
rect -1791 -527 -1761 -505
rect -1695 -527 -1665 -505
rect -1599 -527 -1569 -505
rect -1503 -527 -1473 -505
rect -1407 -527 -1377 -505
rect -1311 -527 -1281 -505
rect -1215 -527 -1185 -505
rect -1119 -527 -1089 -505
rect -1023 -527 -993 -505
rect -927 -527 -897 -505
rect -831 -527 -801 -505
rect -735 -527 -705 -505
rect -639 -527 -609 -505
rect -543 -527 -513 -505
rect -447 -527 -417 -505
rect -351 -527 -321 -505
rect -255 -527 -225 -505
rect -159 -527 -129 -505
rect -63 -527 -33 -505
rect 33 -527 63 -505
rect 129 -527 159 -505
rect 225 -527 255 -505
rect 321 -527 351 -505
rect 417 -527 447 -505
rect 513 -527 543 -505
rect 609 -527 639 -505
rect 705 -527 735 -505
rect 801 -527 831 -505
rect 897 -527 927 -505
rect 993 -527 1023 -505
rect 1089 -527 1119 -505
rect 1185 -527 1215 -505
rect 1281 -527 1311 -505
rect 1377 -527 1407 -505
rect 1473 -527 1503 -505
rect 1569 -527 1599 -505
rect 1665 -527 1695 -505
rect 1761 -527 1791 -505
rect 1857 -527 1887 -505
rect -1887 -749 -1857 -727
rect -1791 -749 -1761 -727
rect -1695 -749 -1665 -727
rect -1599 -749 -1569 -727
rect -1503 -749 -1473 -727
rect -1407 -749 -1377 -727
rect -1311 -749 -1281 -727
rect -1215 -749 -1185 -727
rect -1119 -749 -1089 -727
rect -1023 -749 -993 -727
rect -927 -749 -897 -727
rect -831 -749 -801 -727
rect -735 -749 -705 -727
rect -639 -749 -609 -727
rect -543 -749 -513 -727
rect -447 -749 -417 -727
rect -351 -749 -321 -727
rect -255 -749 -225 -727
rect -159 -749 -129 -727
rect -63 -749 -33 -727
rect 33 -749 63 -727
rect 129 -749 159 -727
rect 225 -749 255 -727
rect 321 -749 351 -727
rect 417 -749 447 -727
rect 513 -749 543 -727
rect 609 -749 639 -727
rect 705 -749 735 -727
rect 801 -749 831 -727
rect 897 -749 927 -727
rect 993 -749 1023 -727
rect 1089 -749 1119 -727
rect 1185 -749 1215 -727
rect 1281 -749 1311 -727
rect 1377 -749 1407 -727
rect 1473 -749 1503 -727
rect 1569 -749 1599 -727
rect 1665 -749 1695 -727
rect 1761 -749 1791 -727
rect 1857 -753 1887 -727
<< locali >>
rect -2051 867 -1955 901
rect 1955 867 2051 901
rect 2017 805 2051 867
rect -1937 715 -1903 731
rect -1937 523 -1903 539
rect -1841 715 -1807 731
rect -1841 523 -1807 539
rect -1745 715 -1711 731
rect -1745 523 -1711 539
rect -1649 715 -1615 731
rect -1649 523 -1615 539
rect -1553 715 -1519 731
rect -1553 523 -1519 539
rect -1457 715 -1423 731
rect -1457 523 -1423 539
rect -1361 715 -1327 731
rect -1361 523 -1327 539
rect -1265 715 -1231 731
rect -1265 523 -1231 539
rect -1169 715 -1135 731
rect -1169 523 -1135 539
rect -1073 715 -1039 731
rect -1073 523 -1039 539
rect -977 715 -943 731
rect -977 523 -943 539
rect -881 715 -847 731
rect -881 523 -847 539
rect -785 715 -751 731
rect -785 523 -751 539
rect -689 715 -655 731
rect -689 523 -655 539
rect -593 715 -559 731
rect -593 523 -559 539
rect -497 715 -463 731
rect -497 523 -463 539
rect -401 715 -367 731
rect -401 523 -367 539
rect -305 715 -271 731
rect -305 523 -271 539
rect -209 715 -175 731
rect -209 523 -175 539
rect -113 715 -79 731
rect -113 523 -79 539
rect -17 715 17 731
rect -17 523 17 539
rect 79 715 113 731
rect 79 523 113 539
rect 175 715 209 731
rect 175 523 209 539
rect 271 715 305 731
rect 271 523 305 539
rect 367 715 401 731
rect 367 523 401 539
rect 463 715 497 731
rect 463 523 497 539
rect 559 715 593 731
rect 559 523 593 539
rect 655 715 689 731
rect 655 523 689 539
rect 751 715 785 731
rect 751 523 785 539
rect 847 715 881 731
rect 847 523 881 539
rect 943 715 977 731
rect 943 523 977 539
rect 1039 715 1073 731
rect 1039 523 1073 539
rect 1135 715 1169 731
rect 1135 523 1169 539
rect 1231 715 1265 731
rect 1231 523 1265 539
rect 1327 715 1361 731
rect 1327 523 1361 539
rect 1423 715 1457 731
rect 1423 523 1457 539
rect 1519 715 1553 731
rect 1519 523 1553 539
rect 1615 715 1649 731
rect 1615 523 1649 539
rect 1711 715 1745 731
rect 1711 523 1745 539
rect 1807 715 1841 731
rect 1807 523 1841 539
rect 1903 715 1937 731
rect 1903 523 1937 539
rect -1937 297 -1903 313
rect -1937 105 -1903 121
rect -1841 297 -1807 313
rect -1841 105 -1807 121
rect -1745 297 -1711 313
rect -1745 105 -1711 121
rect -1649 297 -1615 313
rect -1649 105 -1615 121
rect -1553 297 -1519 313
rect -1553 105 -1519 121
rect -1457 297 -1423 313
rect -1457 105 -1423 121
rect -1361 297 -1327 313
rect -1361 105 -1327 121
rect -1265 297 -1231 313
rect -1265 105 -1231 121
rect -1169 297 -1135 313
rect -1169 105 -1135 121
rect -1073 297 -1039 313
rect -1073 105 -1039 121
rect -977 297 -943 313
rect -977 105 -943 121
rect -881 297 -847 313
rect -881 105 -847 121
rect -785 297 -751 313
rect -785 105 -751 121
rect -689 297 -655 313
rect -689 105 -655 121
rect -593 297 -559 313
rect -593 105 -559 121
rect -497 297 -463 313
rect -497 105 -463 121
rect -401 297 -367 313
rect -401 105 -367 121
rect -305 297 -271 313
rect -305 105 -271 121
rect -209 297 -175 313
rect -209 105 -175 121
rect -113 297 -79 313
rect -113 105 -79 121
rect -17 297 17 313
rect -17 105 17 121
rect 79 297 113 313
rect 79 105 113 121
rect 175 297 209 313
rect 175 105 209 121
rect 271 297 305 313
rect 271 105 305 121
rect 367 297 401 313
rect 367 105 401 121
rect 463 297 497 313
rect 463 105 497 121
rect 559 297 593 313
rect 559 105 593 121
rect 655 297 689 313
rect 655 105 689 121
rect 751 297 785 313
rect 751 105 785 121
rect 847 297 881 313
rect 847 105 881 121
rect 943 297 977 313
rect 943 105 977 121
rect 1039 297 1073 313
rect 1039 105 1073 121
rect 1135 297 1169 313
rect 1135 105 1169 121
rect 1231 297 1265 313
rect 1231 105 1265 121
rect 1327 297 1361 313
rect 1327 105 1361 121
rect 1423 297 1457 313
rect 1423 105 1457 121
rect 1519 297 1553 313
rect 1519 105 1553 121
rect 1615 297 1649 313
rect 1615 105 1649 121
rect 1711 297 1745 313
rect 1711 105 1745 121
rect 1807 297 1841 313
rect 1807 105 1841 121
rect 1903 297 1937 313
rect 1903 105 1937 121
rect -1937 -121 -1903 -105
rect -1937 -313 -1903 -297
rect -1841 -121 -1807 -105
rect -1841 -313 -1807 -297
rect -1745 -121 -1711 -105
rect -1745 -313 -1711 -297
rect -1649 -121 -1615 -105
rect -1649 -313 -1615 -297
rect -1553 -121 -1519 -105
rect -1553 -313 -1519 -297
rect -1457 -121 -1423 -105
rect -1457 -313 -1423 -297
rect -1361 -121 -1327 -105
rect -1361 -313 -1327 -297
rect -1265 -121 -1231 -105
rect -1265 -313 -1231 -297
rect -1169 -121 -1135 -105
rect -1169 -313 -1135 -297
rect -1073 -121 -1039 -105
rect -1073 -313 -1039 -297
rect -977 -121 -943 -105
rect -977 -313 -943 -297
rect -881 -121 -847 -105
rect -881 -313 -847 -297
rect -785 -121 -751 -105
rect -785 -313 -751 -297
rect -689 -121 -655 -105
rect -689 -313 -655 -297
rect -593 -121 -559 -105
rect -593 -313 -559 -297
rect -497 -121 -463 -105
rect -497 -313 -463 -297
rect -401 -121 -367 -105
rect -401 -313 -367 -297
rect -305 -121 -271 -105
rect -305 -313 -271 -297
rect -209 -121 -175 -105
rect -209 -313 -175 -297
rect -113 -121 -79 -105
rect -113 -313 -79 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 79 -121 113 -105
rect 79 -313 113 -297
rect 175 -121 209 -105
rect 175 -313 209 -297
rect 271 -121 305 -105
rect 271 -313 305 -297
rect 367 -121 401 -105
rect 367 -313 401 -297
rect 463 -121 497 -105
rect 463 -313 497 -297
rect 559 -121 593 -105
rect 559 -313 593 -297
rect 655 -121 689 -105
rect 655 -313 689 -297
rect 751 -121 785 -105
rect 751 -313 785 -297
rect 847 -121 881 -105
rect 847 -313 881 -297
rect 943 -121 977 -105
rect 943 -313 977 -297
rect 1039 -121 1073 -105
rect 1039 -313 1073 -297
rect 1135 -121 1169 -105
rect 1135 -313 1169 -297
rect 1231 -121 1265 -105
rect 1231 -313 1265 -297
rect 1327 -121 1361 -105
rect 1327 -313 1361 -297
rect 1423 -121 1457 -105
rect 1423 -313 1457 -297
rect 1519 -121 1553 -105
rect 1519 -313 1553 -297
rect 1615 -121 1649 -105
rect 1615 -313 1649 -297
rect 1711 -121 1745 -105
rect 1711 -313 1745 -297
rect 1807 -121 1841 -105
rect 1807 -313 1841 -297
rect 1903 -121 1937 -105
rect 1903 -313 1937 -297
rect -1937 -539 -1903 -523
rect -1937 -731 -1903 -715
rect -1841 -539 -1807 -523
rect -1841 -731 -1807 -715
rect -1745 -539 -1711 -523
rect -1745 -731 -1711 -715
rect -1649 -539 -1615 -523
rect -1649 -731 -1615 -715
rect -1553 -539 -1519 -523
rect -1553 -731 -1519 -715
rect -1457 -539 -1423 -523
rect -1457 -731 -1423 -715
rect -1361 -539 -1327 -523
rect -1361 -731 -1327 -715
rect -1265 -539 -1231 -523
rect -1265 -731 -1231 -715
rect -1169 -539 -1135 -523
rect -1169 -731 -1135 -715
rect -1073 -539 -1039 -523
rect -1073 -731 -1039 -715
rect -977 -539 -943 -523
rect -977 -731 -943 -715
rect -881 -539 -847 -523
rect -881 -731 -847 -715
rect -785 -539 -751 -523
rect -785 -731 -751 -715
rect -689 -539 -655 -523
rect -689 -731 -655 -715
rect -593 -539 -559 -523
rect -593 -731 -559 -715
rect -497 -539 -463 -523
rect -497 -731 -463 -715
rect -401 -539 -367 -523
rect -401 -731 -367 -715
rect -305 -539 -271 -523
rect -305 -731 -271 -715
rect -209 -539 -175 -523
rect -209 -731 -175 -715
rect -113 -539 -79 -523
rect -113 -731 -79 -715
rect -17 -539 17 -523
rect -17 -731 17 -715
rect 79 -539 113 -523
rect 79 -731 113 -715
rect 175 -539 209 -523
rect 175 -731 209 -715
rect 271 -539 305 -523
rect 271 -731 305 -715
rect 367 -539 401 -523
rect 367 -731 401 -715
rect 463 -539 497 -523
rect 463 -731 497 -715
rect 559 -539 593 -523
rect 559 -731 593 -715
rect 655 -539 689 -523
rect 655 -731 689 -715
rect 751 -539 785 -523
rect 751 -731 785 -715
rect 847 -539 881 -523
rect 847 -731 881 -715
rect 943 -539 977 -523
rect 943 -731 977 -715
rect 1039 -539 1073 -523
rect 1039 -731 1073 -715
rect 1135 -539 1169 -523
rect 1135 -731 1169 -715
rect 1231 -539 1265 -523
rect 1231 -731 1265 -715
rect 1327 -539 1361 -523
rect 1327 -731 1361 -715
rect 1423 -539 1457 -523
rect 1423 -731 1457 -715
rect 1519 -539 1553 -523
rect 1519 -731 1553 -715
rect 1615 -539 1649 -523
rect 1615 -731 1649 -715
rect 1711 -539 1745 -523
rect 1711 -731 1745 -715
rect 1807 -539 1841 -523
rect 1807 -731 1841 -715
rect 1903 -539 1937 -523
rect 1903 -731 1937 -715
rect 2017 -867 2051 -805
rect -2051 -901 -1955 -867
rect 1955 -901 2051 -867
<< viali >>
rect -1937 539 -1903 715
rect -1841 539 -1807 715
rect -1745 539 -1711 715
rect -1649 539 -1615 715
rect -1553 539 -1519 715
rect -1457 539 -1423 715
rect -1361 539 -1327 715
rect -1265 539 -1231 715
rect -1169 539 -1135 715
rect -1073 539 -1039 715
rect -977 539 -943 715
rect -881 539 -847 715
rect -785 539 -751 715
rect -689 539 -655 715
rect -593 539 -559 715
rect -497 539 -463 715
rect -401 539 -367 715
rect -305 539 -271 715
rect -209 539 -175 715
rect -113 539 -79 715
rect -17 539 17 715
rect 79 539 113 715
rect 175 539 209 715
rect 271 539 305 715
rect 367 539 401 715
rect 463 539 497 715
rect 559 539 593 715
rect 655 539 689 715
rect 751 539 785 715
rect 847 539 881 715
rect 943 539 977 715
rect 1039 539 1073 715
rect 1135 539 1169 715
rect 1231 539 1265 715
rect 1327 539 1361 715
rect 1423 539 1457 715
rect 1519 539 1553 715
rect 1615 539 1649 715
rect 1711 539 1745 715
rect 1807 539 1841 715
rect 1903 539 1937 715
rect -1937 121 -1903 297
rect -1841 121 -1807 297
rect -1745 121 -1711 297
rect -1649 121 -1615 297
rect -1553 121 -1519 297
rect -1457 121 -1423 297
rect -1361 121 -1327 297
rect -1265 121 -1231 297
rect -1169 121 -1135 297
rect -1073 121 -1039 297
rect -977 121 -943 297
rect -881 121 -847 297
rect -785 121 -751 297
rect -689 121 -655 297
rect -593 121 -559 297
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect 559 121 593 297
rect 655 121 689 297
rect 751 121 785 297
rect 847 121 881 297
rect 943 121 977 297
rect 1039 121 1073 297
rect 1135 121 1169 297
rect 1231 121 1265 297
rect 1327 121 1361 297
rect 1423 121 1457 297
rect 1519 121 1553 297
rect 1615 121 1649 297
rect 1711 121 1745 297
rect 1807 121 1841 297
rect 1903 121 1937 297
rect -1937 -297 -1903 -121
rect -1841 -297 -1807 -121
rect -1745 -297 -1711 -121
rect -1649 -297 -1615 -121
rect -1553 -297 -1519 -121
rect -1457 -297 -1423 -121
rect -1361 -297 -1327 -121
rect -1265 -297 -1231 -121
rect -1169 -297 -1135 -121
rect -1073 -297 -1039 -121
rect -977 -297 -943 -121
rect -881 -297 -847 -121
rect -785 -297 -751 -121
rect -689 -297 -655 -121
rect -593 -297 -559 -121
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect 559 -297 593 -121
rect 655 -297 689 -121
rect 751 -297 785 -121
rect 847 -297 881 -121
rect 943 -297 977 -121
rect 1039 -297 1073 -121
rect 1135 -297 1169 -121
rect 1231 -297 1265 -121
rect 1327 -297 1361 -121
rect 1423 -297 1457 -121
rect 1519 -297 1553 -121
rect 1615 -297 1649 -121
rect 1711 -297 1745 -121
rect 1807 -297 1841 -121
rect 1903 -297 1937 -121
rect -1937 -715 -1903 -539
rect -1841 -715 -1807 -539
rect -1745 -715 -1711 -539
rect -1649 -715 -1615 -539
rect -1553 -715 -1519 -539
rect -1457 -715 -1423 -539
rect -1361 -715 -1327 -539
rect -1265 -715 -1231 -539
rect -1169 -715 -1135 -539
rect -1073 -715 -1039 -539
rect -977 -715 -943 -539
rect -881 -715 -847 -539
rect -785 -715 -751 -539
rect -689 -715 -655 -539
rect -593 -715 -559 -539
rect -497 -715 -463 -539
rect -401 -715 -367 -539
rect -305 -715 -271 -539
rect -209 -715 -175 -539
rect -113 -715 -79 -539
rect -17 -715 17 -539
rect 79 -715 113 -539
rect 175 -715 209 -539
rect 271 -715 305 -539
rect 367 -715 401 -539
rect 463 -715 497 -539
rect 559 -715 593 -539
rect 655 -715 689 -539
rect 751 -715 785 -539
rect 847 -715 881 -539
rect 943 -715 977 -539
rect 1039 -715 1073 -539
rect 1135 -715 1169 -539
rect 1231 -715 1265 -539
rect 1327 -715 1361 -539
rect 1423 -715 1457 -539
rect 1519 -715 1553 -539
rect 1615 -715 1649 -539
rect 1711 -715 1745 -539
rect 1807 -715 1841 -539
rect 1903 -715 1937 -539
<< metal1 >>
rect -1943 715 -1897 727
rect -1943 539 -1937 715
rect -1903 539 -1897 715
rect -1943 527 -1897 539
rect -1847 715 -1801 727
rect -1847 539 -1841 715
rect -1807 539 -1801 715
rect -1847 527 -1801 539
rect -1751 715 -1705 727
rect -1751 539 -1745 715
rect -1711 539 -1705 715
rect -1751 527 -1705 539
rect -1655 715 -1609 727
rect -1655 539 -1649 715
rect -1615 539 -1609 715
rect -1655 527 -1609 539
rect -1559 715 -1513 727
rect -1559 539 -1553 715
rect -1519 539 -1513 715
rect -1559 527 -1513 539
rect -1463 715 -1417 727
rect -1463 539 -1457 715
rect -1423 539 -1417 715
rect -1463 527 -1417 539
rect -1367 715 -1321 727
rect -1367 539 -1361 715
rect -1327 539 -1321 715
rect -1367 527 -1321 539
rect -1271 715 -1225 727
rect -1271 539 -1265 715
rect -1231 539 -1225 715
rect -1271 527 -1225 539
rect -1175 715 -1129 727
rect -1175 539 -1169 715
rect -1135 539 -1129 715
rect -1175 527 -1129 539
rect -1079 715 -1033 727
rect -1079 539 -1073 715
rect -1039 539 -1033 715
rect -1079 527 -1033 539
rect -983 715 -937 727
rect -983 539 -977 715
rect -943 539 -937 715
rect -983 527 -937 539
rect -887 715 -841 727
rect -887 539 -881 715
rect -847 539 -841 715
rect -887 527 -841 539
rect -791 715 -745 727
rect -791 539 -785 715
rect -751 539 -745 715
rect -791 527 -745 539
rect -695 715 -649 727
rect -695 539 -689 715
rect -655 539 -649 715
rect -695 527 -649 539
rect -599 715 -553 727
rect -599 539 -593 715
rect -559 539 -553 715
rect -599 527 -553 539
rect -503 715 -457 727
rect -503 539 -497 715
rect -463 539 -457 715
rect -503 527 -457 539
rect -407 715 -361 727
rect -407 539 -401 715
rect -367 539 -361 715
rect -407 527 -361 539
rect -311 715 -265 727
rect -311 539 -305 715
rect -271 539 -265 715
rect -311 527 -265 539
rect -215 715 -169 727
rect -215 539 -209 715
rect -175 539 -169 715
rect -215 527 -169 539
rect -119 715 -73 727
rect -119 539 -113 715
rect -79 539 -73 715
rect -119 527 -73 539
rect -23 715 23 727
rect -23 539 -17 715
rect 17 539 23 715
rect -23 527 23 539
rect 73 715 119 727
rect 73 539 79 715
rect 113 539 119 715
rect 73 527 119 539
rect 169 715 215 727
rect 169 539 175 715
rect 209 539 215 715
rect 169 527 215 539
rect 265 715 311 727
rect 265 539 271 715
rect 305 539 311 715
rect 265 527 311 539
rect 361 715 407 727
rect 361 539 367 715
rect 401 539 407 715
rect 361 527 407 539
rect 457 715 503 727
rect 457 539 463 715
rect 497 539 503 715
rect 457 527 503 539
rect 553 715 599 727
rect 553 539 559 715
rect 593 539 599 715
rect 553 527 599 539
rect 649 715 695 727
rect 649 539 655 715
rect 689 539 695 715
rect 649 527 695 539
rect 745 715 791 727
rect 745 539 751 715
rect 785 539 791 715
rect 745 527 791 539
rect 841 715 887 727
rect 841 539 847 715
rect 881 539 887 715
rect 841 527 887 539
rect 937 715 983 727
rect 937 539 943 715
rect 977 539 983 715
rect 937 527 983 539
rect 1033 715 1079 727
rect 1033 539 1039 715
rect 1073 539 1079 715
rect 1033 527 1079 539
rect 1129 715 1175 727
rect 1129 539 1135 715
rect 1169 539 1175 715
rect 1129 527 1175 539
rect 1225 715 1271 727
rect 1225 539 1231 715
rect 1265 539 1271 715
rect 1225 527 1271 539
rect 1321 715 1367 727
rect 1321 539 1327 715
rect 1361 539 1367 715
rect 1321 527 1367 539
rect 1417 715 1463 727
rect 1417 539 1423 715
rect 1457 539 1463 715
rect 1417 527 1463 539
rect 1513 715 1559 727
rect 1513 539 1519 715
rect 1553 539 1559 715
rect 1513 527 1559 539
rect 1609 715 1655 727
rect 1609 539 1615 715
rect 1649 539 1655 715
rect 1609 527 1655 539
rect 1705 715 1751 727
rect 1705 539 1711 715
rect 1745 539 1751 715
rect 1705 527 1751 539
rect 1801 715 1847 727
rect 1801 539 1807 715
rect 1841 539 1847 715
rect 1801 527 1847 539
rect 1897 715 1943 727
rect 1897 539 1903 715
rect 1937 539 1943 715
rect 1897 527 1943 539
rect -1943 297 -1897 309
rect -1943 121 -1937 297
rect -1903 121 -1897 297
rect -1943 109 -1897 121
rect -1847 297 -1801 309
rect -1847 121 -1841 297
rect -1807 121 -1801 297
rect -1847 109 -1801 121
rect -1751 297 -1705 309
rect -1751 121 -1745 297
rect -1711 121 -1705 297
rect -1751 109 -1705 121
rect -1655 297 -1609 309
rect -1655 121 -1649 297
rect -1615 121 -1609 297
rect -1655 109 -1609 121
rect -1559 297 -1513 309
rect -1559 121 -1553 297
rect -1519 121 -1513 297
rect -1559 109 -1513 121
rect -1463 297 -1417 309
rect -1463 121 -1457 297
rect -1423 121 -1417 297
rect -1463 109 -1417 121
rect -1367 297 -1321 309
rect -1367 121 -1361 297
rect -1327 121 -1321 297
rect -1367 109 -1321 121
rect -1271 297 -1225 309
rect -1271 121 -1265 297
rect -1231 121 -1225 297
rect -1271 109 -1225 121
rect -1175 297 -1129 309
rect -1175 121 -1169 297
rect -1135 121 -1129 297
rect -1175 109 -1129 121
rect -1079 297 -1033 309
rect -1079 121 -1073 297
rect -1039 121 -1033 297
rect -1079 109 -1033 121
rect -983 297 -937 309
rect -983 121 -977 297
rect -943 121 -937 297
rect -983 109 -937 121
rect -887 297 -841 309
rect -887 121 -881 297
rect -847 121 -841 297
rect -887 109 -841 121
rect -791 297 -745 309
rect -791 121 -785 297
rect -751 121 -745 297
rect -791 109 -745 121
rect -695 297 -649 309
rect -695 121 -689 297
rect -655 121 -649 297
rect -695 109 -649 121
rect -599 297 -553 309
rect -599 121 -593 297
rect -559 121 -553 297
rect -599 109 -553 121
rect -503 297 -457 309
rect -503 121 -497 297
rect -463 121 -457 297
rect -503 109 -457 121
rect -407 297 -361 309
rect -407 121 -401 297
rect -367 121 -361 297
rect -407 109 -361 121
rect -311 297 -265 309
rect -311 121 -305 297
rect -271 121 -265 297
rect -311 109 -265 121
rect -215 297 -169 309
rect -215 121 -209 297
rect -175 121 -169 297
rect -215 109 -169 121
rect -119 297 -73 309
rect -119 121 -113 297
rect -79 121 -73 297
rect -119 109 -73 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 73 297 119 309
rect 73 121 79 297
rect 113 121 119 297
rect 73 109 119 121
rect 169 297 215 309
rect 169 121 175 297
rect 209 121 215 297
rect 169 109 215 121
rect 265 297 311 309
rect 265 121 271 297
rect 305 121 311 297
rect 265 109 311 121
rect 361 297 407 309
rect 361 121 367 297
rect 401 121 407 297
rect 361 109 407 121
rect 457 297 503 309
rect 457 121 463 297
rect 497 121 503 297
rect 457 109 503 121
rect 553 297 599 309
rect 553 121 559 297
rect 593 121 599 297
rect 553 109 599 121
rect 649 297 695 309
rect 649 121 655 297
rect 689 121 695 297
rect 649 109 695 121
rect 745 297 791 309
rect 745 121 751 297
rect 785 121 791 297
rect 745 109 791 121
rect 841 297 887 309
rect 841 121 847 297
rect 881 121 887 297
rect 841 109 887 121
rect 937 297 983 309
rect 937 121 943 297
rect 977 121 983 297
rect 937 109 983 121
rect 1033 297 1079 309
rect 1033 121 1039 297
rect 1073 121 1079 297
rect 1033 109 1079 121
rect 1129 297 1175 309
rect 1129 121 1135 297
rect 1169 121 1175 297
rect 1129 109 1175 121
rect 1225 297 1271 309
rect 1225 121 1231 297
rect 1265 121 1271 297
rect 1225 109 1271 121
rect 1321 297 1367 309
rect 1321 121 1327 297
rect 1361 121 1367 297
rect 1321 109 1367 121
rect 1417 297 1463 309
rect 1417 121 1423 297
rect 1457 121 1463 297
rect 1417 109 1463 121
rect 1513 297 1559 309
rect 1513 121 1519 297
rect 1553 121 1559 297
rect 1513 109 1559 121
rect 1609 297 1655 309
rect 1609 121 1615 297
rect 1649 121 1655 297
rect 1609 109 1655 121
rect 1705 297 1751 309
rect 1705 121 1711 297
rect 1745 121 1751 297
rect 1705 109 1751 121
rect 1801 297 1847 309
rect 1801 121 1807 297
rect 1841 121 1847 297
rect 1801 109 1847 121
rect 1897 297 1943 309
rect 1897 121 1903 297
rect 1937 121 1943 297
rect 1897 109 1943 121
rect -1943 -121 -1897 -109
rect -1943 -297 -1937 -121
rect -1903 -297 -1897 -121
rect -1943 -309 -1897 -297
rect -1847 -121 -1801 -109
rect -1847 -297 -1841 -121
rect -1807 -297 -1801 -121
rect -1847 -309 -1801 -297
rect -1751 -121 -1705 -109
rect -1751 -297 -1745 -121
rect -1711 -297 -1705 -121
rect -1751 -309 -1705 -297
rect -1655 -121 -1609 -109
rect -1655 -297 -1649 -121
rect -1615 -297 -1609 -121
rect -1655 -309 -1609 -297
rect -1559 -121 -1513 -109
rect -1559 -297 -1553 -121
rect -1519 -297 -1513 -121
rect -1559 -309 -1513 -297
rect -1463 -121 -1417 -109
rect -1463 -297 -1457 -121
rect -1423 -297 -1417 -121
rect -1463 -309 -1417 -297
rect -1367 -121 -1321 -109
rect -1367 -297 -1361 -121
rect -1327 -297 -1321 -121
rect -1367 -309 -1321 -297
rect -1271 -121 -1225 -109
rect -1271 -297 -1265 -121
rect -1231 -297 -1225 -121
rect -1271 -309 -1225 -297
rect -1175 -121 -1129 -109
rect -1175 -297 -1169 -121
rect -1135 -297 -1129 -121
rect -1175 -309 -1129 -297
rect -1079 -121 -1033 -109
rect -1079 -297 -1073 -121
rect -1039 -297 -1033 -121
rect -1079 -309 -1033 -297
rect -983 -121 -937 -109
rect -983 -297 -977 -121
rect -943 -297 -937 -121
rect -983 -309 -937 -297
rect -887 -121 -841 -109
rect -887 -297 -881 -121
rect -847 -297 -841 -121
rect -887 -309 -841 -297
rect -791 -121 -745 -109
rect -791 -297 -785 -121
rect -751 -297 -745 -121
rect -791 -309 -745 -297
rect -695 -121 -649 -109
rect -695 -297 -689 -121
rect -655 -297 -649 -121
rect -695 -309 -649 -297
rect -599 -121 -553 -109
rect -599 -297 -593 -121
rect -559 -297 -553 -121
rect -599 -309 -553 -297
rect -503 -121 -457 -109
rect -503 -297 -497 -121
rect -463 -297 -457 -121
rect -503 -309 -457 -297
rect -407 -121 -361 -109
rect -407 -297 -401 -121
rect -367 -297 -361 -121
rect -407 -309 -361 -297
rect -311 -121 -265 -109
rect -311 -297 -305 -121
rect -271 -297 -265 -121
rect -311 -309 -265 -297
rect -215 -121 -169 -109
rect -215 -297 -209 -121
rect -175 -297 -169 -121
rect -215 -309 -169 -297
rect -119 -121 -73 -109
rect -119 -297 -113 -121
rect -79 -297 -73 -121
rect -119 -309 -73 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 73 -121 119 -109
rect 73 -297 79 -121
rect 113 -297 119 -121
rect 73 -309 119 -297
rect 169 -121 215 -109
rect 169 -297 175 -121
rect 209 -297 215 -121
rect 169 -309 215 -297
rect 265 -121 311 -109
rect 265 -297 271 -121
rect 305 -297 311 -121
rect 265 -309 311 -297
rect 361 -121 407 -109
rect 361 -297 367 -121
rect 401 -297 407 -121
rect 361 -309 407 -297
rect 457 -121 503 -109
rect 457 -297 463 -121
rect 497 -297 503 -121
rect 457 -309 503 -297
rect 553 -121 599 -109
rect 553 -297 559 -121
rect 593 -297 599 -121
rect 553 -309 599 -297
rect 649 -121 695 -109
rect 649 -297 655 -121
rect 689 -297 695 -121
rect 649 -309 695 -297
rect 745 -121 791 -109
rect 745 -297 751 -121
rect 785 -297 791 -121
rect 745 -309 791 -297
rect 841 -121 887 -109
rect 841 -297 847 -121
rect 881 -297 887 -121
rect 841 -309 887 -297
rect 937 -121 983 -109
rect 937 -297 943 -121
rect 977 -297 983 -121
rect 937 -309 983 -297
rect 1033 -121 1079 -109
rect 1033 -297 1039 -121
rect 1073 -297 1079 -121
rect 1033 -309 1079 -297
rect 1129 -121 1175 -109
rect 1129 -297 1135 -121
rect 1169 -297 1175 -121
rect 1129 -309 1175 -297
rect 1225 -121 1271 -109
rect 1225 -297 1231 -121
rect 1265 -297 1271 -121
rect 1225 -309 1271 -297
rect 1321 -121 1367 -109
rect 1321 -297 1327 -121
rect 1361 -297 1367 -121
rect 1321 -309 1367 -297
rect 1417 -121 1463 -109
rect 1417 -297 1423 -121
rect 1457 -297 1463 -121
rect 1417 -309 1463 -297
rect 1513 -121 1559 -109
rect 1513 -297 1519 -121
rect 1553 -297 1559 -121
rect 1513 -309 1559 -297
rect 1609 -121 1655 -109
rect 1609 -297 1615 -121
rect 1649 -297 1655 -121
rect 1609 -309 1655 -297
rect 1705 -121 1751 -109
rect 1705 -297 1711 -121
rect 1745 -297 1751 -121
rect 1705 -309 1751 -297
rect 1801 -121 1847 -109
rect 1801 -297 1807 -121
rect 1841 -297 1847 -121
rect 1801 -309 1847 -297
rect 1897 -121 1943 -109
rect 1897 -297 1903 -121
rect 1937 -297 1943 -121
rect 1897 -309 1943 -297
rect -1943 -539 -1897 -527
rect -1943 -715 -1937 -539
rect -1903 -715 -1897 -539
rect -1943 -727 -1897 -715
rect -1847 -539 -1801 -527
rect -1847 -715 -1841 -539
rect -1807 -715 -1801 -539
rect -1847 -727 -1801 -715
rect -1751 -539 -1705 -527
rect -1751 -715 -1745 -539
rect -1711 -715 -1705 -539
rect -1751 -727 -1705 -715
rect -1655 -539 -1609 -527
rect -1655 -715 -1649 -539
rect -1615 -715 -1609 -539
rect -1655 -727 -1609 -715
rect -1559 -539 -1513 -527
rect -1559 -715 -1553 -539
rect -1519 -715 -1513 -539
rect -1559 -727 -1513 -715
rect -1463 -539 -1417 -527
rect -1463 -715 -1457 -539
rect -1423 -715 -1417 -539
rect -1463 -727 -1417 -715
rect -1367 -539 -1321 -527
rect -1367 -715 -1361 -539
rect -1327 -715 -1321 -539
rect -1367 -727 -1321 -715
rect -1271 -539 -1225 -527
rect -1271 -715 -1265 -539
rect -1231 -715 -1225 -539
rect -1271 -727 -1225 -715
rect -1175 -539 -1129 -527
rect -1175 -715 -1169 -539
rect -1135 -715 -1129 -539
rect -1175 -727 -1129 -715
rect -1079 -539 -1033 -527
rect -1079 -715 -1073 -539
rect -1039 -715 -1033 -539
rect -1079 -727 -1033 -715
rect -983 -539 -937 -527
rect -983 -715 -977 -539
rect -943 -715 -937 -539
rect -983 -727 -937 -715
rect -887 -539 -841 -527
rect -887 -715 -881 -539
rect -847 -715 -841 -539
rect -887 -727 -841 -715
rect -791 -539 -745 -527
rect -791 -715 -785 -539
rect -751 -715 -745 -539
rect -791 -727 -745 -715
rect -695 -539 -649 -527
rect -695 -715 -689 -539
rect -655 -715 -649 -539
rect -695 -727 -649 -715
rect -599 -539 -553 -527
rect -599 -715 -593 -539
rect -559 -715 -553 -539
rect -599 -727 -553 -715
rect -503 -539 -457 -527
rect -503 -715 -497 -539
rect -463 -715 -457 -539
rect -503 -727 -457 -715
rect -407 -539 -361 -527
rect -407 -715 -401 -539
rect -367 -715 -361 -539
rect -407 -727 -361 -715
rect -311 -539 -265 -527
rect -311 -715 -305 -539
rect -271 -715 -265 -539
rect -311 -727 -265 -715
rect -215 -539 -169 -527
rect -215 -715 -209 -539
rect -175 -715 -169 -539
rect -215 -727 -169 -715
rect -119 -539 -73 -527
rect -119 -715 -113 -539
rect -79 -715 -73 -539
rect -119 -727 -73 -715
rect -23 -539 23 -527
rect -23 -715 -17 -539
rect 17 -715 23 -539
rect -23 -727 23 -715
rect 73 -539 119 -527
rect 73 -715 79 -539
rect 113 -715 119 -539
rect 73 -727 119 -715
rect 169 -539 215 -527
rect 169 -715 175 -539
rect 209 -715 215 -539
rect 169 -727 215 -715
rect 265 -539 311 -527
rect 265 -715 271 -539
rect 305 -715 311 -539
rect 265 -727 311 -715
rect 361 -539 407 -527
rect 361 -715 367 -539
rect 401 -715 407 -539
rect 361 -727 407 -715
rect 457 -539 503 -527
rect 457 -715 463 -539
rect 497 -715 503 -539
rect 457 -727 503 -715
rect 553 -539 599 -527
rect 553 -715 559 -539
rect 593 -715 599 -539
rect 553 -727 599 -715
rect 649 -539 695 -527
rect 649 -715 655 -539
rect 689 -715 695 -539
rect 649 -727 695 -715
rect 745 -539 791 -527
rect 745 -715 751 -539
rect 785 -715 791 -539
rect 745 -727 791 -715
rect 841 -539 887 -527
rect 841 -715 847 -539
rect 881 -715 887 -539
rect 841 -727 887 -715
rect 937 -539 983 -527
rect 937 -715 943 -539
rect 977 -715 983 -539
rect 937 -727 983 -715
rect 1033 -539 1079 -527
rect 1033 -715 1039 -539
rect 1073 -715 1079 -539
rect 1033 -727 1079 -715
rect 1129 -539 1175 -527
rect 1129 -715 1135 -539
rect 1169 -715 1175 -539
rect 1129 -727 1175 -715
rect 1225 -539 1271 -527
rect 1225 -715 1231 -539
rect 1265 -715 1271 -539
rect 1225 -727 1271 -715
rect 1321 -539 1367 -527
rect 1321 -715 1327 -539
rect 1361 -715 1367 -539
rect 1321 -727 1367 -715
rect 1417 -539 1463 -527
rect 1417 -715 1423 -539
rect 1457 -715 1463 -539
rect 1417 -727 1463 -715
rect 1513 -539 1559 -527
rect 1513 -715 1519 -539
rect 1553 -715 1559 -539
rect 1513 -727 1559 -715
rect 1609 -539 1655 -527
rect 1609 -715 1615 -539
rect 1649 -715 1655 -539
rect 1609 -727 1655 -715
rect 1705 -539 1751 -527
rect 1705 -715 1711 -539
rect 1745 -715 1751 -539
rect 1705 -727 1751 -715
rect 1801 -539 1847 -527
rect 1801 -715 1807 -539
rect 1841 -715 1847 -539
rect 1801 -727 1847 -715
rect 1897 -539 1943 -527
rect 1897 -715 1903 -539
rect 1937 -715 1943 -539
rect 1897 -727 1943 -715
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -2034 -884 2034 884
string parameters w 1 l 0.150 m 4 nf 40 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
