magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect -211 -309 211 309
<< pmos >>
rect -15 -90 15 90
<< pdiff >>
rect -73 78 -15 90
rect -73 -78 -61 78
rect -27 -78 -15 78
rect -73 -90 -15 -78
rect 15 78 73 90
rect 15 -78 27 78
rect 61 -78 73 78
rect 15 -90 73 -78
<< pdiffc >>
rect -61 -78 -27 78
rect 27 -78 61 78
<< nsubdiff >>
rect -141 239 -79 273
rect 79 239 175 273
rect 141 177 175 239
rect 141 -239 175 -177
<< nsubdiffcont >>
rect -79 239 79 273
rect 141 -177 175 177
<< poly >>
rect -15 90 15 121
rect -15 -121 15 -90
rect -51 -187 15 -121
<< locali >>
rect -141 239 -79 273
rect 79 239 175 273
rect 141 177 175 239
rect -61 78 -27 94
rect -61 -94 -27 -78
rect 27 78 61 94
rect 27 -94 61 -78
rect 141 -239 175 -177
<< viali >>
rect -61 -78 -27 78
rect 27 -78 61 78
<< metal1 >>
rect -67 78 -21 90
rect -67 -78 -61 78
rect -27 -78 -21 78
rect -67 -90 -21 -78
rect 21 78 67 90
rect 21 -78 27 78
rect 61 -78 67 78
rect 21 -90 67 -78
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -158 -256 158 256
string parameters w 0.9 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
