magic
tech sky130A
magscale 1 2
timestamp 1623427962
<< nwell >>
rect -263 -303 263 303
<< pmos >>
rect -63 -84 -33 84
rect 33 -84 63 84
<< pdiff >>
rect -125 72 -63 84
rect -125 -72 -113 72
rect -79 -72 -63 72
rect -125 -84 -63 -72
rect -33 72 33 84
rect -33 -72 -17 72
rect 17 -72 33 72
rect -33 -84 33 -72
rect 63 72 125 84
rect 63 -72 79 72
rect 113 -72 125 72
rect 63 -84 125 -72
<< pdiffc >>
rect -113 -72 -79 72
rect -17 -72 17 72
rect 79 -72 113 72
<< nsubdiff >>
rect -227 233 -131 267
rect 131 233 227 267
rect -227 171 -193 233
rect 193 171 227 233
rect -227 -233 -193 -171
rect 193 -233 227 -171
<< nsubdiffcont >>
rect -131 233 131 267
rect -227 -171 -193 171
rect 193 -171 227 171
<< poly >>
rect -63 84 -33 110
rect 33 84 63 110
rect -63 -110 -33 -84
rect 33 -110 63 -84
<< locali >>
rect -227 233 -131 267
rect 131 233 227 267
rect -227 171 -193 233
rect 193 171 227 233
rect -113 72 -79 88
rect -113 -88 -79 -72
rect -17 72 17 88
rect -17 -88 17 -72
rect 79 72 113 88
rect 79 -88 113 -72
rect -227 -233 -193 -171
rect 193 -233 227 -171
<< viali >>
rect -113 -72 -79 72
rect -17 -72 17 72
rect 79 -72 113 72
<< metal1 >>
rect -119 72 -73 84
rect -119 -72 -113 72
rect -79 -72 -73 72
rect -119 -84 -73 -72
rect -23 72 23 84
rect -23 -72 -17 72
rect 17 -72 23 72
rect -23 -84 23 -72
rect 73 72 119 84
rect 73 -72 79 72
rect 113 -72 119 72
rect 73 -84 119 -72
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -210 -250 210 250
string parameters w 0.84 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
