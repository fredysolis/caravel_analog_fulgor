magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< nwell >>
rect -33 2264 526 2352
rect -33 2261 525 2264
rect -33 2137 307 2261
rect -33 1900 340 2137
rect -33 1576 526 1900
rect -33 -1 526 60
rect -33 -628 0 -1
rect -33 -716 526 -628
<< pwell >>
rect -33 1030 0 1576
rect -33 967 503 1030
rect -33 669 526 967
rect -33 668 503 669
rect -33 60 0 668
<< psubdiff >>
rect 36 1506 434 1540
rect 36 563 70 1027
rect 453 1002 555 1036
rect 424 600 633 634
rect 36 130 70 182
rect 36 96 613 130
<< nsubdiff >>
rect 107 2282 131 2316
rect 393 2282 417 2316
rect 108 -680 132 -646
rect 394 -680 418 -646
<< nsubdiffcont >>
rect 131 2282 393 2316
rect 132 -680 394 -646
<< poly >>
rect 99 1807 230 1824
rect 99 1773 124 1807
rect 192 1773 230 1807
rect 99 1758 230 1773
rect 296 -137 427 -122
rect 296 -171 334 -137
rect 402 -171 427 -137
rect 296 -188 427 -171
<< polycont >>
rect 124 1773 192 1807
rect 334 -171 402 -137
<< locali >>
rect 108 1773 124 1807
rect 192 1773 208 1807
rect 70 1506 434 1540
rect 70 96 434 130
rect 318 -171 334 -137
rect 402 -171 418 -137
<< viali >>
rect 36 2282 131 2316
rect 131 2282 393 2316
rect 393 2282 490 2316
rect 36 2194 490 2228
rect 124 1773 192 1807
rect 36 1036 70 1540
rect 36 1002 555 1036
rect 36 634 70 1002
rect 36 600 1077 634
rect 36 96 70 600
rect 434 96 1112 130
rect 334 -171 402 -137
rect 36 -592 490 -558
rect 36 -680 132 -646
rect 132 -680 394 -646
rect 394 -680 490 -646
<< metal1 >>
rect -33 2316 526 2322
rect -33 2282 36 2316
rect 490 2282 526 2316
rect -33 2228 526 2282
rect -33 2194 36 2228
rect 490 2194 526 2228
rect -33 2188 526 2194
rect 144 2045 190 2188
rect 336 2045 382 2188
rect 102 1761 112 1813
rect 194 1761 204 1813
rect 240 1651 286 1901
rect 30 1540 76 1552
rect 227 1547 237 1651
rect 289 1547 299 1651
rect 30 982 36 1540
rect 70 1042 76 1540
rect 240 1366 286 1547
rect 198 1104 328 1138
rect 70 1036 567 1042
rect 555 1002 567 1036
rect -33 654 36 982
rect 30 96 36 654
rect 70 996 567 1002
rect 70 640 76 996
rect 70 634 1089 640
rect 1077 600 1089 634
rect 70 594 1089 600
rect 70 96 76 594
rect 198 498 328 532
rect 766 519 812 594
rect 958 519 1004 594
rect 657 392 667 511
rect 657 280 667 346
rect 719 280 729 511
rect 849 281 859 512
rect 911 281 921 512
rect 30 84 76 96
rect 240 89 286 270
rect 714 192 954 232
rect 422 130 1124 136
rect 422 96 434 130
rect 1112 96 1124 130
rect 422 90 1124 96
rect 227 -15 237 89
rect 289 -15 299 89
rect 240 -219 286 -15
rect 322 -177 332 -125
rect 414 -177 424 -125
rect 144 -552 190 -408
rect 336 -552 382 -399
rect -33 -558 526 -552
rect -33 -592 36 -558
rect 490 -592 526 -558
rect -33 -646 526 -592
rect -33 -680 36 -646
rect 490 -680 526 -646
rect -33 -686 526 -680
<< via1 >>
rect 112 1807 194 1813
rect 112 1773 124 1807
rect 124 1773 192 1807
rect 192 1773 194 1807
rect 112 1761 194 1773
rect 237 1547 289 1651
rect 667 280 719 511
rect 859 281 911 512
rect 237 -15 289 89
rect 332 -137 414 -125
rect 332 -171 334 -137
rect 334 -171 402 -137
rect 402 -171 414 -137
rect 332 -177 414 -171
<< metal2 >>
rect 102 1814 214 1824
rect 102 1748 214 1758
rect 237 1651 289 1661
rect 340 1653 396 1663
rect 289 1570 340 1629
rect 237 1537 289 1547
rect 396 1570 398 1629
rect 340 1532 396 1542
rect 497 1323 553 1333
rect 359 1239 497 1299
rect 497 1201 553 1211
rect 667 511 719 521
rect 859 512 911 522
rect 470 396 582 404
rect 360 394 667 396
rect 360 338 470 394
rect 582 338 667 394
rect 360 336 667 338
rect 470 328 582 336
rect 719 281 859 511
rect 719 280 911 281
rect 667 270 719 280
rect 859 271 911 280
rect 130 94 186 104
rect 128 7 130 66
rect 237 89 289 99
rect 186 7 237 66
rect 130 -26 186 -17
rect 237 -25 289 -15
rect 312 -122 424 -112
rect 312 -188 424 -178
<< via2 >>
rect 102 1813 214 1814
rect 102 1761 112 1813
rect 112 1761 194 1813
rect 194 1761 214 1813
rect 102 1758 214 1761
rect 340 1542 396 1653
rect 497 1211 553 1323
rect 470 338 582 394
rect 130 -17 186 94
rect 312 -125 424 -122
rect 312 -177 332 -125
rect 332 -177 414 -125
rect 414 -177 424 -125
rect 312 -178 424 -177
<< metal3 >>
rect 92 1814 224 1819
rect 92 1758 102 1814
rect 214 1758 224 1814
rect 92 1753 224 1758
rect 128 99 188 1753
rect 330 1653 406 1658
rect 330 1542 340 1653
rect 396 1542 406 1653
rect 330 1537 406 1542
rect 120 94 196 99
rect 120 -17 130 94
rect 186 -17 196 94
rect 120 -22 196 -17
rect 338 -117 398 1537
rect 495 1328 555 1333
rect 487 1323 563 1328
rect 487 1211 497 1323
rect 553 1211 563 1323
rect 487 1206 563 1211
rect 495 399 555 1206
rect 460 394 592 399
rect 460 338 470 394
rect 582 338 592 394
rect 460 333 592 338
rect 495 323 555 333
rect 302 -122 434 -117
rect 302 -178 312 -122
rect 424 -178 434 -122
rect 302 -183 434 -178
use sky130_fd_pr__nfet_01v8_2BS854  sky130_fd_pr__nfet_01v8_2BS854_0
timestamp 1624049879
transform 1 0 836 0 1 395
box -311 -335 311 335
use sky130_fd_pr__pfet_01v8_MJG8BZ  sky130_fd_pr__pfet_01v8_MJG8BZ_0
timestamp 1624049879
transform 1 0 263 0 1 1950
box -263 -314 263 314
use sky130_fd_pr__pfet_01v8_MJG8BZ  sky130_fd_pr__pfet_01v8_MJG8BZ_1
timestamp 1624049879
transform -1 0 263 0 -1 -314
box -263 -314 263 314
use sky130_fd_pr__nfet_01v8_KU9PSX  sky130_fd_pr__nfet_01v8_KU9PSX_1
timestamp 1624049879
transform 1 0 263 0 1 1271
box -263 -305 263 305
use sky130_fd_pr__nfet_01v8_KU9PSX  sky130_fd_pr__nfet_01v8_KU9PSX_0
timestamp 1624049879
transform 1 0 263 0 -1 365
box -263 -305 263 305
<< labels >>
rlabel metal1 -33 654 36 982 1 vss
rlabel metal1 -33 2228 526 2282 1 vdd
rlabel metal3 128 94 188 1758 1 Q
rlabel metal3 338 -122 398 1542 1 nQ
rlabel metal1 198 1104 328 1138 1 D
rlabel metal1 198 498 328 532 1 nD
rlabel metal1 -33 -646 526 -592 1 vdd
rlabel metal1 714 192 954 232 1 CLK
<< end >>
