* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_1_MACBVW VSUBS m3_n2650_n13200# m3_n7969_n2600# m3_7988_8000#
+ m3_2669_n7900# m3_n13288_n2600# m3_n2650_2700# m3_2669_2700# m3_n13288_n13200# m3_n7969_n13200#
+ m3_n13288_8000# m3_7988_2700# m3_n2650_n7900# m3_7988_n7900# m3_2669_n13200# m3_n7969_8000#
+ m3_n13288_2700# m3_n7969_n7900# m3_n13288_n7900# m3_2669_n2600# m3_n7969_2700# m3_7988_n13200#
+ c1_n13188_n13100# m3_7988_n2600# m3_n2650_n2600# m3_n2650_8000# m3_2669_8000#
X0 c1_n13188_n13100# m3_2669_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X1 c1_n13188_n13100# m3_n2650_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X2 c1_n13188_n13100# m3_2669_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X3 c1_n13188_n13100# m3_n13288_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X4 c1_n13188_n13100# m3_n7969_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X5 c1_n13188_n13100# m3_n13288_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X6 c1_n13188_n13100# m3_2669_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X7 c1_n13188_n13100# m3_7988_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X8 c1_n13188_n13100# m3_2669_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X9 c1_n13188_n13100# m3_7988_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X10 c1_n13188_n13100# m3_n7969_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X11 c1_n13188_n13100# m3_7988_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X12 c1_n13188_n13100# m3_n7969_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X13 c1_n13188_n13100# m3_7988_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X14 c1_n13188_n13100# m3_n13288_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X15 c1_n13188_n13100# m3_n7969_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X16 c1_n13188_n13100# m3_n2650_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X17 c1_n13188_n13100# m3_n2650_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X18 c1_n13188_n13100# m3_n2650_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X19 c1_n13188_n13100# m3_7988_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X20 c1_n13188_n13100# m3_n13288_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X21 c1_n13188_n13100# m3_n13288_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X22 c1_n13188_n13100# m3_n7969_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X23 c1_n13188_n13100# m3_n2650_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X24 c1_n13188_n13100# m3_2669_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
C0 m3_n7969_n2600# c1_n13188_n13100# 58.86fF
C1 m3_7988_n2600# m3_7988_n7900# 3.39fF
C2 m3_2669_n7900# m3_7988_n7900# 2.73fF
C3 m3_2669_2700# m3_7988_2700# 2.73fF
C4 m3_n7969_n7900# m3_n2650_n7900# 2.73fF
C5 m3_7988_8000# m3_7988_2700# 3.39fF
C6 c1_n13188_n13100# m3_n2650_n7900# 58.86fF
C7 m3_n7969_8000# m3_n7969_2700# 3.28fF
C8 m3_2669_8000# m3_n2650_8000# 2.73fF
C9 m3_n13288_8000# m3_n7969_8000# 2.73fF
C10 m3_2669_8000# c1_n13188_n13100# 58.61fF
C11 m3_n13288_n13200# c1_n13188_n13100# 58.36fF
C12 m3_7988_n13200# m3_7988_n7900# 3.39fF
C13 m3_n7969_n2600# m3_n7969_2700# 3.28fF
C14 m3_2669_n7900# m3_n2650_n7900# 2.73fF
C15 m3_n2650_8000# m3_n2650_2700# 3.28fF
C16 m3_n2650_n13200# m3_n2650_n7900# 3.28fF
C17 m3_n13288_n13200# m3_n7969_n13200# 2.73fF
C18 m3_n13288_2700# m3_n13288_n2600# 3.28fF
C19 c1_n13188_n13100# m3_n2650_2700# 58.86fF
C20 m3_n7969_n2600# m3_n2650_n2600# 2.73fF
C21 m3_n13288_2700# c1_n13188_n13100# 58.61fF
C22 m3_n13288_n13200# m3_n13288_n7900# 3.28fF
C23 m3_n2650_8000# c1_n13188_n13100# 58.61fF
C24 m3_2669_n13200# c1_n13188_n13100# 58.61fF
C25 c1_n13188_n13100# m3_2669_n2600# 58.86fF
C26 c1_n13188_n13100# m3_n13288_n2600# 58.61fF
C27 m3_n7969_n7900# c1_n13188_n13100# 58.86fF
C28 m3_n2650_n2600# m3_n2650_n7900# 3.28fF
C29 m3_n7969_n7900# m3_n7969_n13200# 3.28fF
C30 c1_n13188_n13100# m3_n7969_n13200# 58.61fF
C31 m3_2669_n2600# m3_7988_n2600# 2.73fF
C32 c1_n13188_n13100# m3_7988_2700# 61.01fF
C33 m3_2669_n7900# m3_2669_n13200# 3.28fF
C34 m3_2669_8000# m3_2669_2700# 3.28fF
C35 m3_n13288_n7900# m3_n13288_n2600# 3.28fF
C36 m3_2669_n7900# m3_2669_n2600# 3.28fF
C37 m3_7988_8000# m3_2669_8000# 2.73fF
C38 c1_n13188_n13100# m3_7988_n2600# 61.01fF
C39 m3_n7969_2700# m3_n2650_2700# 2.73fF
C40 m3_n7969_n7900# m3_n13288_n7900# 2.73fF
C41 m3_n2650_n13200# m3_2669_n13200# 2.73fF
C42 c1_n13188_n13100# m3_n13288_n7900# 58.61fF
C43 m3_n13288_2700# m3_n7969_2700# 2.73fF
C44 m3_2669_n7900# c1_n13188_n13100# 58.86fF
C45 m3_n2650_n13200# c1_n13188_n13100# 58.61fF
C46 m3_n7969_8000# m3_n2650_8000# 2.73fF
C47 m3_n13288_8000# m3_n13288_2700# 3.28fF
C48 c1_n13188_n13100# m3_n7969_2700# 58.86fF
C49 m3_7988_n2600# m3_7988_2700# 3.39fF
C50 c1_n13188_n13100# m3_7988_n7900# 61.01fF
C51 m3_2669_2700# m3_n2650_2700# 2.73fF
C52 m3_n2650_n2600# m3_n2650_2700# 3.28fF
C53 m3_n7969_8000# c1_n13188_n13100# 58.61fF
C54 m3_n13288_8000# c1_n13188_n13100# 58.36fF
C55 m3_n2650_n13200# m3_n7969_n13200# 2.73fF
C56 m3_2669_2700# m3_2669_n2600# 3.28fF
C57 m3_n2650_n2600# m3_2669_n2600# 2.73fF
C58 m3_7988_n13200# m3_2669_n13200# 2.73fF
C59 m3_2669_2700# c1_n13188_n13100# 58.86fF
C60 m3_n2650_n2600# c1_n13188_n13100# 58.86fF
C61 m3_n7969_n2600# m3_n13288_n2600# 2.73fF
C62 m3_7988_8000# c1_n13188_n13100# 60.75fF
C63 m3_7988_n13200# c1_n13188_n13100# 60.75fF
C64 m3_n7969_n2600# m3_n7969_n7900# 3.28fF
C65 c1_n13188_n13100# VSUBS 2.51fF
C66 m3_7988_n13200# VSUBS 12.57fF
C67 m3_2669_n13200# VSUBS 12.37fF
C68 m3_n2650_n13200# VSUBS 12.37fF
C69 m3_n7969_n13200# VSUBS 12.37fF
C70 m3_n13288_n13200# VSUBS 12.37fF
C71 m3_7988_n7900# VSUBS 12.57fF
C72 m3_2669_n7900# VSUBS 12.37fF
C73 m3_n2650_n7900# VSUBS 12.37fF
C74 m3_n7969_n7900# VSUBS 12.37fF
C75 m3_n13288_n7900# VSUBS 12.37fF
C76 m3_7988_n2600# VSUBS 12.57fF
C77 m3_2669_n2600# VSUBS 12.37fF
C78 m3_n2650_n2600# VSUBS 12.37fF
C79 m3_n7969_n2600# VSUBS 12.37fF
C80 m3_n13288_n2600# VSUBS 12.37fF
C81 m3_7988_2700# VSUBS 12.57fF
C82 m3_2669_2700# VSUBS 12.37fF
C83 m3_n2650_2700# VSUBS 12.37fF
C84 m3_n7969_2700# VSUBS 12.37fF
C85 m3_n13288_2700# VSUBS 12.37fF
C86 m3_7988_8000# VSUBS 12.57fF
C87 m3_2669_8000# VSUBS 12.37fF
C88 m3_n2650_8000# VSUBS 12.37fF
C89 m3_n7969_8000# VSUBS 12.37fF
C90 m3_n13288_8000# VSUBS 12.37fF
.ends

.subckt cap1_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_MACBVW_0 VSUBS out out out out out out out out out out
+ out out out out out out out out out out out in out out out out sky130_fd_pr__cap_mim_m3_1_MACBVW
C0 in out 2.17fF
C1 in VSUBS -10.03fF
C2 out VSUBS 62.40fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_W3JTNJ VSUBS m3_n6469_n2100# c1_n6369_n6300# m3_2169_n6400#
+ m3_n2150_n6400# c1_2269_n6300# m3_n6469_2200# m3_n2150_n2100# c1_n2050_n6300# m3_n2150_2200#
+ m3_n6469_n6400#
X0 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2 c1_n2050_n6300# m3_n2150_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 c1_n6369_n6300# m3_n6469_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X4 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X5 c1_n6369_n6300# m3_n6469_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X6 c1_n2050_n6300# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X7 c1_n2050_n6300# m3_n2150_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X8 c1_n6369_n6300# m3_n6469_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
C0 m3_n2150_n6400# c1_n2050_n6300# 38.10fF
C1 m3_n2150_2200# c1_n2050_n6300# 38.10fF
C2 c1_n6369_n6300# c1_n2050_n6300# 1.99fF
C3 c1_2269_n6300# c1_n2050_n6300# 1.99fF
C4 m3_2169_n6400# m3_n2150_n6400# 1.75fF
C5 m3_2169_n6400# m3_n2150_2200# 1.75fF
C6 m3_2169_n6400# c1_2269_n6300# 121.67fF
C7 m3_n6469_n2100# m3_n6469_2200# 2.63fF
C8 m3_n6469_n2100# m3_n6469_n6400# 2.63fF
C9 m3_n6469_n2100# m3_n2150_n2100# 1.75fF
C10 m3_n2150_n2100# c1_n2050_n6300# 38.10fF
C11 m3_2169_n6400# m3_n2150_n2100# 1.75fF
C12 m3_n6469_2200# m3_n2150_2200# 1.75fF
C13 m3_n6469_n6400# m3_n2150_n6400# 1.75fF
C14 m3_n2150_n2100# m3_n2150_n6400# 2.63fF
C15 m3_n6469_2200# c1_n6369_n6300# 38.10fF
C16 m3_n2150_2200# m3_n2150_n2100# 2.63fF
C17 m3_n6469_n6400# c1_n6369_n6300# 38.10fF
C18 m3_n6469_n2100# c1_n6369_n6300# 38.10fF
C19 c1_2269_n6300# VSUBS 0.16fF
C20 c1_n2050_n6300# VSUBS 0.16fF
C21 c1_n6369_n6300# VSUBS 0.16fF
C22 m3_n2150_n6400# VSUBS 8.68fF
C23 m3_n6469_n6400# VSUBS 8.68fF
C24 m3_n2150_n2100# VSUBS 8.68fF
C25 m3_n6469_n2100# VSUBS 8.68fF
C26 m3_2169_n6400# VSUBS 26.86fF
C27 m3_n2150_2200# VSUBS 8.68fF
C28 m3_n6469_2200# VSUBS 8.68fF
.ends

.subckt cap2_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_W3JTNJ_0 VSUBS out in out out in out out in out out sky130_fd_pr__cap_mim_m3_1_W3JTNJ
C0 out in 8.08fF
C1 in VSUBS -16.59fF
C2 out VSUBS 13.00fF
.ends

.subckt sky130_fd_pr__res_high_po_5p73_X44RQA a_n573_2292# w_n739_n2890# a_n573_n2724#
X0 a_n573_n2724# a_n573_2292# w_n739_n2890# sky130_fd_pr__res_high_po_5p73 l=2.292e+07u
C0 a_n573_n2724# w_n739_n2890# 1.98fF
C1 a_n573_2292# w_n739_n2890# 1.98fF
.ends

.subckt res_loop_filter vss out in
Xsky130_fd_pr__res_high_po_5p73_X44RQA_0 in vss out sky130_fd_pr__res_high_po_5p73_X44RQA
C0 out vss 3.87fF
C1 in vss 3.02fF
.ends

.subckt loop_filter vc_pex in vss
Xcap1_loop_filter_0 vss vc_pex vss cap1_loop_filter
Xcap2_loop_filter_0 vss in vss cap2_loop_filter
Xres_loop_filter_0 vss res_loop_filter_2/out in res_loop_filter
Xres_loop_filter_1 vss res_loop_filter_2/out vc_pex res_loop_filter
Xres_loop_filter_2 vss res_loop_filter_2/out vc_pex res_loop_filter
C0 in vc_pex 0.18fF
C1 vc_pex vss -38.13fF
C2 res_loop_filter_2/out vss 8.49fF
C3 in vss -18.79fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4ML9WA VSUBS a_429_n486# w_n2457_n634# a_887_n486#
+ a_n29_n486# a_1345_n486# a_n2261_n512# a_1803_n486# a_n487_n486# a_n945_n486# a_n2319_n486#
+ a_n1403_n486# a_2261_n486# a_n1861_n486#
X0 a_2261_n486# a_n2261_n512# a_1803_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X1 a_n945_n486# a_n2261_n512# a_n1403_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X2 a_429_n486# a_n2261_n512# a_n29_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X3 a_1803_n486# a_n2261_n512# a_1345_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X4 a_887_n486# a_n2261_n512# a_429_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X5 a_n487_n486# a_n2261_n512# a_n945_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X6 a_n1403_n486# a_n2261_n512# a_n1861_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X7 a_n1861_n486# a_n2261_n512# a_n2319_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X8 a_n29_n486# a_n2261_n512# a_n487_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X9 a_1345_n486# a_n2261_n512# a_887_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
C0 w_n2457_n634# a_n1403_n486# 0.02fF
C1 w_n2457_n634# a_1345_n486# 0.02fF
C2 w_n2457_n634# a_n1861_n486# 0.02fF
C3 w_n2457_n634# a_2261_n486# 0.02fF
C4 w_n2457_n634# a_1803_n486# 0.02fF
C5 w_n2457_n634# a_n2319_n486# 0.02fF
C6 w_n2457_n634# a_n945_n486# 0.02fF
C7 w_n2457_n634# a_n487_n486# 0.02fF
C8 w_n2457_n634# a_887_n486# 0.02fF
C9 w_n2457_n634# a_429_n486# 0.02fF
C10 w_n2457_n634# a_n29_n486# 0.02fF
C11 a_2261_n486# VSUBS 0.03fF
C12 a_1803_n486# VSUBS 0.03fF
C13 a_1345_n486# VSUBS 0.03fF
C14 a_887_n486# VSUBS 0.03fF
C15 a_429_n486# VSUBS 0.03fF
C16 a_n29_n486# VSUBS 0.03fF
C17 a_n487_n486# VSUBS 0.03fF
C18 a_n945_n486# VSUBS 0.03fF
C19 a_n1403_n486# VSUBS 0.03fF
C20 a_n1861_n486# VSUBS 0.03fF
C21 a_n2319_n486# VSUBS 0.03fF
C22 a_n2261_n512# VSUBS 4.27fF
C23 w_n2457_n634# VSUBS 21.34fF
.ends

.subckt sky130_fd_pr__nfet_01v8_YCGG98 a_n1041_n75# a_n561_n75# a_1167_n75# a_303_n75#
+ a_687_n75# a_n849_n75# a_n369_n75# a_975_n75# a_111_n75# a_495_n75# a_n1137_n75#
+ a_n657_n75# a_n177_n75# a_783_n75# a_n945_n75# a_n465_n75# a_207_n75# a_1071_n75#
+ a_591_n75# a_15_n75# a_n753_n75# w_n1367_n285# a_n273_n75# a_879_n75# a_399_n75#
+ a_n1229_n75# a_n81_n75# a_n1167_n101#
X0 a_207_n75# a_n1167_n101# a_111_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_303_n75# a_n1167_n101# a_207_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_399_n75# a_n1167_n101# a_303_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_495_n75# a_n1167_n101# a_399_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_591_n75# a_n1167_n101# a_495_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_783_n75# a_n1167_n101# a_687_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_687_n75# a_n1167_n101# a_591_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_879_n75# a_n1167_n101# a_783_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_975_n75# a_n1167_n101# a_879_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_n1041_n75# a_n1167_n101# a_n1137_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_n1137_n75# a_n1167_n101# a_n1229_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n561_n75# a_n1167_n101# a_n657_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_1071_n75# a_n1167_n101# a_975_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n945_n75# a_n1167_n101# a_n1041_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n753_n75# a_n1167_n101# a_n849_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n657_n75# a_n1167_n101# a_n753_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n465_n75# a_n1167_n101# a_n561_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n369_n75# a_n1167_n101# a_n465_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_1167_n75# a_n1167_n101# a_1071_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n849_n75# a_n1167_n101# a_n945_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X20 a_15_n75# a_n1167_n101# a_n81_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X21 a_n81_n75# a_n1167_n101# a_n177_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X22 a_111_n75# a_n1167_n101# a_15_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X23 a_n273_n75# a_n1167_n101# a_n369_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X24 a_n177_n75# a_n1167_n101# a_n273_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
C0 a_303_n75# a_207_n75# 0.22fF
C1 a_n945_n75# a_n657_n75# 0.05fF
C2 a_15_n75# a_n177_n75# 0.08fF
C3 a_n465_n75# a_n657_n75# 0.08fF
C4 a_n1041_n75# a_n657_n75# 0.03fF
C5 a_n369_n75# a_n177_n75# 0.08fF
C6 a_n465_n75# a_n273_n75# 0.08fF
C7 a_n945_n75# a_n753_n75# 0.08fF
C8 a_111_n75# a_n273_n75# 0.03fF
C9 a_n1137_n75# a_n945_n75# 0.08fF
C10 a_n465_n75# a_n753_n75# 0.05fF
C11 a_n1041_n75# a_n753_n75# 0.05fF
C12 a_n81_n75# a_n273_n75# 0.08fF
C13 a_783_n75# a_975_n75# 0.08fF
C14 a_879_n75# a_1167_n75# 0.05fF
C15 a_n1041_n75# a_n1137_n75# 0.22fF
C16 a_495_n75# a_303_n75# 0.08fF
C17 a_111_n75# a_303_n75# 0.08fF
C18 a_n849_n75# a_n945_n75# 0.22fF
C19 a_1071_n75# a_975_n75# 0.22fF
C20 a_n81_n75# a_303_n75# 0.03fF
C21 a_n849_n75# a_n465_n75# 0.03fF
C22 a_n849_n75# a_n1041_n75# 0.08fF
C23 a_687_n75# a_303_n75# 0.03fF
C24 a_n561_n75# a_n369_n75# 0.08fF
C25 a_1071_n75# a_783_n75# 0.05fF
C26 a_n273_n75# a_n177_n75# 0.22fF
C27 a_495_n75# a_207_n75# 0.05fF
C28 a_111_n75# a_207_n75# 0.22fF
C29 a_687_n75# a_975_n75# 0.05fF
C30 a_n81_n75# a_207_n75# 0.05fF
C31 a_495_n75# a_783_n75# 0.05fF
C32 a_687_n75# a_783_n75# 0.22fF
C33 a_591_n75# a_399_n75# 0.08fF
C34 a_n1041_n75# a_n945_n75# 0.22fF
C35 a_15_n75# a_399_n75# 0.03fF
C36 a_n561_n75# a_n657_n75# 0.22fF
C37 a_879_n75# a_591_n75# 0.05fF
C38 a_687_n75# a_1071_n75# 0.03fF
C39 a_n561_n75# a_n273_n75# 0.05fF
C40 a_15_n75# a_n369_n75# 0.03fF
C41 a_495_n75# a_111_n75# 0.03fF
C42 a_n561_n75# a_n753_n75# 0.08fF
C43 a_207_n75# a_n177_n75# 0.03fF
C44 a_n81_n75# a_n465_n75# 0.03fF
C45 a_111_n75# a_n81_n75# 0.08fF
C46 a_687_n75# a_495_n75# 0.08fF
C47 a_n849_n75# a_n561_n75# 0.05fF
C48 a_1167_n75# a_975_n75# 0.08fF
C49 a_n465_n75# a_n177_n75# 0.05fF
C50 a_111_n75# a_n177_n75# 0.05fF
C51 a_1167_n75# a_783_n75# 0.03fF
C52 a_n81_n75# a_n177_n75# 0.22fF
C53 a_n369_n75# a_n657_n75# 0.05fF
C54 a_15_n75# a_n273_n75# 0.05fF
C55 a_303_n75# a_399_n75# 0.22fF
C56 a_1071_n75# a_1167_n75# 0.22fF
C57 a_n369_n75# a_n273_n75# 0.22fF
C58 a_n369_n75# a_n753_n75# 0.03fF
C59 a_n561_n75# a_n945_n75# 0.03fF
C60 a_591_n75# a_303_n75# 0.05fF
C61 a_15_n75# a_303_n75# 0.05fF
C62 a_n561_n75# a_n465_n75# 0.22fF
C63 a_n1137_n75# a_n1229_n75# 0.22fF
C64 a_207_n75# a_399_n75# 0.08fF
C65 a_879_n75# a_975_n75# 0.22fF
C66 a_n849_n75# a_n1229_n75# 0.03fF
C67 a_783_n75# a_399_n75# 0.03fF
C68 a_591_n75# a_975_n75# 0.03fF
C69 a_591_n75# a_207_n75# 0.03fF
C70 a_879_n75# a_783_n75# 0.22fF
C71 a_15_n75# a_207_n75# 0.08fF
C72 a_n657_n75# a_n273_n75# 0.03fF
C73 a_783_n75# a_591_n75# 0.08fF
C74 a_1071_n75# a_879_n75# 0.08fF
C75 a_n753_n75# a_n657_n75# 0.22fF
C76 a_n561_n75# a_n177_n75# 0.03fF
C77 a_495_n75# a_399_n75# 0.22fF
C78 a_111_n75# a_399_n75# 0.05fF
C79 a_n945_n75# a_n1229_n75# 0.05fF
C80 a_879_n75# a_495_n75# 0.03fF
C81 a_n849_n75# a_n657_n75# 0.08fF
C82 a_n1137_n75# a_n753_n75# 0.03fF
C83 a_687_n75# a_399_n75# 0.05fF
C84 a_n465_n75# a_n369_n75# 0.22fF
C85 a_495_n75# a_591_n75# 0.22fF
C86 a_111_n75# a_15_n75# 0.22fF
C87 a_n1041_n75# a_n1229_n75# 0.08fF
C88 a_687_n75# a_879_n75# 0.08fF
C89 a_n81_n75# a_15_n75# 0.22fF
C90 a_n849_n75# a_n753_n75# 0.22fF
C91 a_n81_n75# a_n369_n75# 0.05fF
C92 a_687_n75# a_591_n75# 0.22fF
C93 a_n849_n75# a_n1137_n75# 0.05fF
C94 a_1167_n75# w_n1367_n285# 0.10fF
C95 a_1071_n75# w_n1367_n285# 0.07fF
C96 a_975_n75# w_n1367_n285# 0.06fF
C97 a_879_n75# w_n1367_n285# 0.05fF
C98 a_783_n75# w_n1367_n285# 0.04fF
C99 a_687_n75# w_n1367_n285# 0.04fF
C100 a_591_n75# w_n1367_n285# 0.04fF
C101 a_495_n75# w_n1367_n285# 0.04fF
C102 a_399_n75# w_n1367_n285# 0.04fF
C103 a_303_n75# w_n1367_n285# 0.04fF
C104 a_207_n75# w_n1367_n285# 0.04fF
C105 a_111_n75# w_n1367_n285# 0.04fF
C106 a_15_n75# w_n1367_n285# 0.04fF
C107 a_n81_n75# w_n1367_n285# 0.04fF
C108 a_n177_n75# w_n1367_n285# 0.04fF
C109 a_n273_n75# w_n1367_n285# 0.04fF
C110 a_n369_n75# w_n1367_n285# 0.04fF
C111 a_n465_n75# w_n1367_n285# 0.04fF
C112 a_n561_n75# w_n1367_n285# 0.04fF
C113 a_n657_n75# w_n1367_n285# 0.04fF
C114 a_n753_n75# w_n1367_n285# 0.04fF
C115 a_n849_n75# w_n1367_n285# 0.04fF
C116 a_n945_n75# w_n1367_n285# 0.04fF
C117 a_n1041_n75# w_n1367_n285# 0.04fF
C118 a_n1137_n75# w_n1367_n285# 0.04fF
C119 a_n1229_n75# w_n1367_n285# 0.04fF
C120 a_n1167_n101# w_n1367_n285# 2.55fF
.ends

.subckt sky130_fd_pr__nfet_01v8_MUHGM9 a_33_n101# a_n129_n75# a_735_n75# a_255_n75#
+ a_n417_n75# a_n989_n75# a_63_n75# a_543_n75# a_n705_n75# a_n225_n75# a_n33_n75#
+ a_831_n75# a_351_n75# a_n927_n101# a_n513_n75# a_n897_n75# w_n1127_n285# a_639_n75#
+ a_159_n75# a_n801_n75# a_n321_n75# a_927_n75# a_447_n75# a_n609_n75#
X0 a_63_n75# a_33_n101# a_n33_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_927_n75# a_33_n101# a_831_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_n33_n75# a_n927_n101# a_n129_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_159_n75# a_33_n101# a_63_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_255_n75# a_33_n101# a_159_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_351_n75# a_33_n101# a_255_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_447_n75# a_33_n101# a_351_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_543_n75# a_33_n101# a_447_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_735_n75# a_33_n101# a_639_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_831_n75# a_33_n101# a_735_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_639_n75# a_33_n101# a_543_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n321_n75# a_n927_n101# a_n417_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_n801_n75# a_n927_n101# a_n897_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n705_n75# a_n927_n101# a_n801_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n513_n75# a_n927_n101# a_n609_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n417_n75# a_n927_n101# a_n513_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n225_n75# a_n927_n101# a_n321_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n129_n75# a_n927_n101# a_n225_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_n897_n75# a_n927_n101# a_n989_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n609_n75# a_n927_n101# a_n705_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
C0 a_n609_n75# a_n417_n75# 0.08fF
C1 a_n801_n75# a_n513_n75# 0.05fF
C2 a_63_n75# a_n33_n75# 0.22fF
C3 a_351_n75# a_639_n75# 0.05fF
C4 a_n225_n75# a_n417_n75# 0.08fF
C5 a_831_n75# a_639_n75# 0.08fF
C6 a_255_n75# a_639_n75# 0.03fF
C7 a_351_n75# a_543_n75# 0.08fF
C8 a_n129_n75# a_n513_n75# 0.03fF
C9 a_351_n75# a_63_n75# 0.05fF
C10 a_831_n75# a_543_n75# 0.05fF
C11 a_255_n75# a_543_n75# 0.05fF
C12 a_n321_n75# a_n513_n75# 0.08fF
C13 a_n705_n75# a_n609_n75# 0.22fF
C14 a_255_n75# a_63_n75# 0.08fF
C15 a_n989_n75# a_n705_n75# 0.05fF
C16 a_927_n75# a_831_n75# 0.22fF
C17 a_n129_n75# a_63_n75# 0.08fF
C18 a_447_n75# a_351_n75# 0.22fF
C19 a_n801_n75# a_n897_n75# 0.22fF
C20 a_n321_n75# a_63_n75# 0.03fF
C21 a_447_n75# a_831_n75# 0.03fF
C22 a_447_n75# a_255_n75# 0.08fF
C23 a_351_n75# a_n33_n75# 0.03fF
C24 a_n513_n75# a_n417_n75# 0.22fF
C25 a_255_n75# a_n33_n75# 0.05fF
C26 a_n129_n75# a_n33_n75# 0.22fF
C27 a_n321_n75# a_n33_n75# 0.05fF
C28 a_n989_n75# a_n609_n75# 0.03fF
C29 a_n927_n101# a_33_n101# 0.08fF
C30 a_255_n75# a_351_n75# 0.22fF
C31 a_n225_n75# a_n609_n75# 0.03fF
C32 a_735_n75# a_639_n75# 0.22fF
C33 a_n705_n75# a_n513_n75# 0.08fF
C34 a_n129_n75# a_255_n75# 0.03fF
C35 a_n225_n75# a_159_n75# 0.03fF
C36 a_735_n75# a_543_n75# 0.08fF
C37 a_n33_n75# a_n417_n75# 0.03fF
C38 a_n129_n75# a_n321_n75# 0.08fF
C39 a_735_n75# a_927_n75# 0.08fF
C40 a_n801_n75# a_n417_n75# 0.03fF
C41 a_447_n75# a_735_n75# 0.05fF
C42 a_n705_n75# a_n897_n75# 0.08fF
C43 a_n609_n75# a_n513_n75# 0.22fF
C44 a_n129_n75# a_n417_n75# 0.05fF
C45 a_n321_n75# a_n417_n75# 0.22fF
C46 a_n225_n75# a_n513_n75# 0.05fF
C47 a_n801_n75# a_n705_n75# 0.22fF
C48 a_159_n75# a_543_n75# 0.03fF
C49 a_735_n75# a_351_n75# 0.03fF
C50 a_n225_n75# a_63_n75# 0.05fF
C51 a_63_n75# a_159_n75# 0.22fF
C52 a_735_n75# a_831_n75# 0.22fF
C53 a_n897_n75# a_n609_n75# 0.05fF
C54 a_n705_n75# a_n321_n75# 0.03fF
C55 a_n989_n75# a_n897_n75# 0.22fF
C56 a_447_n75# a_159_n75# 0.05fF
C57 a_n225_n75# a_n33_n75# 0.08fF
C58 a_n801_n75# a_n609_n75# 0.08fF
C59 a_159_n75# a_n33_n75# 0.08fF
C60 a_n801_n75# a_n989_n75# 0.08fF
C61 a_543_n75# a_639_n75# 0.22fF
C62 a_n705_n75# a_n417_n75# 0.05fF
C63 a_927_n75# a_639_n75# 0.05fF
C64 a_351_n75# a_159_n75# 0.08fF
C65 a_n321_n75# a_n609_n75# 0.05fF
C66 a_447_n75# a_639_n75# 0.08fF
C67 a_927_n75# a_543_n75# 0.03fF
C68 a_255_n75# a_159_n75# 0.22fF
C69 a_n129_n75# a_n225_n75# 0.22fF
C70 a_n129_n75# a_159_n75# 0.05fF
C71 a_n321_n75# a_n225_n75# 0.22fF
C72 a_447_n75# a_543_n75# 0.22fF
C73 a_n897_n75# a_n513_n75# 0.03fF
C74 a_447_n75# a_63_n75# 0.03fF
C75 a_927_n75# w_n1127_n285# 0.04fF
C76 a_831_n75# w_n1127_n285# 0.04fF
C77 a_735_n75# w_n1127_n285# 0.04fF
C78 a_639_n75# w_n1127_n285# 0.04fF
C79 a_543_n75# w_n1127_n285# 0.04fF
C80 a_447_n75# w_n1127_n285# 0.04fF
C81 a_351_n75# w_n1127_n285# 0.04fF
C82 a_255_n75# w_n1127_n285# 0.04fF
C83 a_159_n75# w_n1127_n285# 0.04fF
C84 a_63_n75# w_n1127_n285# 0.04fF
C85 a_n33_n75# w_n1127_n285# 0.04fF
C86 a_n129_n75# w_n1127_n285# 0.04fF
C87 a_n225_n75# w_n1127_n285# 0.04fF
C88 a_n321_n75# w_n1127_n285# 0.04fF
C89 a_n417_n75# w_n1127_n285# 0.04fF
C90 a_n513_n75# w_n1127_n285# 0.04fF
C91 a_n609_n75# w_n1127_n285# 0.04fF
C92 a_n705_n75# w_n1127_n285# 0.04fF
C93 a_n801_n75# w_n1127_n285# 0.04fF
C94 a_n897_n75# w_n1127_n285# 0.04fF
C95 a_n989_n75# w_n1127_n285# 0.04fF
C96 a_33_n101# w_n1127_n285# 0.99fF
C97 a_n927_n101# w_n1127_n285# 0.99fF
.ends

.subckt sky130_fd_pr__pfet_01v8_NKZXKB VSUBS a_33_n247# a_n801_n150# a_n417_n150#
+ a_351_n150# a_255_n150# a_n705_n150# a_n609_n150# a_159_n150# a_543_n150# a_447_n150#
+ a_831_n150# a_n897_n150# a_n33_n150# a_735_n150# a_n927_n247# a_639_n150# a_n321_n150#
+ a_927_n150# a_n225_n150# a_63_n150# a_n989_n150# a_n513_n150# a_n129_n150# w_n1127_n369#
X0 a_n513_n150# a_n927_n247# a_n609_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_63_n150# a_33_n247# a_n33_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_735_n150# a_33_n247# a_639_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n801_n150# a_n927_n247# a_n897_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n927_n247# a_n225_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n927_n247# a_n513_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_639_n150# a_33_n247# a_543_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n705_n150# a_n927_n247# a_n801_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n33_n150# a_n927_n247# a_n129_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_351_n150# a_33_n247# a_255_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_n609_n150# a_n927_n247# a_n705_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n897_n150# a_n927_n247# a_n989_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_927_n150# a_33_n247# a_831_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_255_n150# a_33_n247# a_159_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n321_n150# a_n927_n247# a_n417_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_543_n150# a_33_n247# a_447_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_831_n150# a_33_n247# a_735_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_159_n150# a_33_n247# a_63_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_n225_n150# a_n927_n247# a_n321_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_447_n150# a_33_n247# a_351_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n705_n150# a_n513_n150# 0.16fF
C1 a_159_n150# a_351_n150# 0.16fF
C2 a_n417_n150# a_n513_n150# 0.43fF
C3 a_n129_n150# a_255_n150# 0.07fF
C4 a_63_n150# a_351_n150# 0.10fF
C5 a_543_n150# a_255_n150# 0.10fF
C6 a_n129_n150# a_n417_n150# 0.10fF
C7 a_447_n150# a_255_n150# 0.16fF
C8 a_n609_n150# a_n705_n150# 0.43fF
C9 a_n225_n150# a_n417_n150# 0.16fF
C10 a_33_n247# a_n927_n247# 0.09fF
C11 a_927_n150# a_639_n150# 0.10fF
C12 a_n609_n150# a_n417_n150# 0.16fF
C13 a_n33_n150# a_n129_n150# 0.43fF
C14 a_735_n150# a_831_n150# 0.43fF
C15 a_n33_n150# a_n225_n150# 0.16fF
C16 a_n129_n150# a_n513_n150# 0.07fF
C17 a_255_n150# a_351_n150# 0.43fF
C18 a_543_n150# a_831_n150# 0.10fF
C19 a_n225_n150# a_n513_n150# 0.10fF
C20 a_n609_n150# a_n513_n150# 0.43fF
C21 a_447_n150# a_831_n150# 0.07fF
C22 a_735_n150# a_543_n150# 0.16fF
C23 a_63_n150# a_159_n150# 0.43fF
C24 a_n225_n150# a_n129_n150# 0.43fF
C25 a_735_n150# a_447_n150# 0.10fF
C26 a_n33_n150# a_351_n150# 0.07fF
C27 a_639_n150# a_255_n150# 0.07fF
C28 a_n609_n150# a_n225_n150# 0.07fF
C29 a_63_n150# a_n321_n150# 0.07fF
C30 a_543_n150# a_447_n150# 0.43fF
C31 a_n897_n150# a_n801_n150# 0.43fF
C32 a_735_n150# a_351_n150# 0.07fF
C33 a_n989_n150# a_n801_n150# 0.16fF
C34 a_n897_n150# a_n989_n150# 0.43fF
C35 a_639_n150# a_831_n150# 0.16fF
C36 a_159_n150# a_255_n150# 0.43fF
C37 a_543_n150# a_351_n150# 0.16fF
C38 a_447_n150# a_351_n150# 0.43fF
C39 a_63_n150# a_255_n150# 0.16fF
C40 a_735_n150# a_639_n150# 0.43fF
C41 a_n321_n150# a_n705_n150# 0.07fF
C42 a_n705_n150# a_n801_n150# 0.43fF
C43 a_n33_n150# a_159_n150# 0.16fF
C44 a_n417_n150# a_n321_n150# 0.43fF
C45 a_n897_n150# a_n705_n150# 0.16fF
C46 a_n417_n150# a_n801_n150# 0.07fF
C47 a_543_n150# a_639_n150# 0.43fF
C48 a_n989_n150# a_n705_n150# 0.10fF
C49 a_n33_n150# a_63_n150# 0.43fF
C50 a_639_n150# a_447_n150# 0.16fF
C51 a_927_n150# a_831_n150# 0.43fF
C52 a_n33_n150# a_n321_n150# 0.10fF
C53 a_n321_n150# a_n513_n150# 0.16fF
C54 a_n801_n150# a_n513_n150# 0.10fF
C55 a_735_n150# a_927_n150# 0.16fF
C56 a_n129_n150# a_159_n150# 0.10fF
C57 a_n897_n150# a_n513_n150# 0.07fF
C58 a_639_n150# a_351_n150# 0.10fF
C59 a_n225_n150# a_159_n150# 0.07fF
C60 a_543_n150# a_159_n150# 0.07fF
C61 a_63_n150# a_n129_n150# 0.16fF
C62 a_n129_n150# a_n321_n150# 0.16fF
C63 a_927_n150# a_543_n150# 0.07fF
C64 a_447_n150# a_159_n150# 0.10fF
C65 a_n417_n150# a_n705_n150# 0.10fF
C66 a_n225_n150# a_63_n150# 0.10fF
C67 a_n33_n150# a_255_n150# 0.10fF
C68 a_n225_n150# a_n321_n150# 0.43fF
C69 a_n609_n150# a_n321_n150# 0.10fF
C70 a_n609_n150# a_n801_n150# 0.16fF
C71 a_447_n150# a_63_n150# 0.07fF
C72 a_n609_n150# a_n897_n150# 0.10fF
C73 a_n33_n150# a_n417_n150# 0.07fF
C74 a_n609_n150# a_n989_n150# 0.07fF
C75 a_927_n150# VSUBS 0.03fF
C76 a_831_n150# VSUBS 0.03fF
C77 a_735_n150# VSUBS 0.03fF
C78 a_639_n150# VSUBS 0.03fF
C79 a_543_n150# VSUBS 0.03fF
C80 a_447_n150# VSUBS 0.03fF
C81 a_351_n150# VSUBS 0.03fF
C82 a_255_n150# VSUBS 0.03fF
C83 a_159_n150# VSUBS 0.03fF
C84 a_63_n150# VSUBS 0.03fF
C85 a_n33_n150# VSUBS 0.03fF
C86 a_n129_n150# VSUBS 0.03fF
C87 a_n225_n150# VSUBS 0.03fF
C88 a_n321_n150# VSUBS 0.03fF
C89 a_n417_n150# VSUBS 0.03fF
C90 a_n513_n150# VSUBS 0.03fF
C91 a_n609_n150# VSUBS 0.03fF
C92 a_n705_n150# VSUBS 0.03fF
C93 a_n801_n150# VSUBS 0.03fF
C94 a_n897_n150# VSUBS 0.03fF
C95 a_n989_n150# VSUBS 0.03fF
C96 a_33_n247# VSUBS 1.04fF
C97 a_n927_n247# VSUBS 1.04fF
C98 w_n1127_n369# VSUBS 6.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_8GRULZ a_n1761_n132# a_1045_n44# a_n1461_n44# a_n1103_n44#
+ a_n29_n44# a_n387_n44# a_1761_n44# a_n1819_n44# a_1403_n44# a_687_n44# w_n1957_n254#
+ a_329_n44# a_n745_n44#
X0 a_329_n44# a_n1761_n132# a_n29_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X1 a_1761_n44# a_n1761_n132# a_1403_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X2 a_n745_n44# a_n1761_n132# a_n1103_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X3 a_1045_n44# a_n1761_n132# a_687_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X4 a_n29_n44# a_n1761_n132# a_n387_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X5 a_n1103_n44# a_n1761_n132# a_n1461_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X6 a_n387_n44# a_n1761_n132# a_n745_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X7 a_687_n44# a_n1761_n132# a_329_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X8 a_1403_n44# a_n1761_n132# a_1045_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X9 a_n1461_n44# a_n1761_n132# a_n1819_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
C0 a_1761_n44# a_1403_n44# 0.04fF
C1 a_n1103_n44# a_n745_n44# 0.04fF
C2 a_1045_n44# a_1403_n44# 0.04fF
C3 a_n387_n44# a_n29_n44# 0.04fF
C4 a_n1103_n44# a_n1461_n44# 0.04fF
C5 a_329_n44# a_687_n44# 0.04fF
C6 a_n1819_n44# a_n1461_n44# 0.04fF
C7 a_n387_n44# a_n745_n44# 0.04fF
C8 a_329_n44# a_n29_n44# 0.04fF
C9 a_1045_n44# a_687_n44# 0.04fF
C10 a_1761_n44# w_n1957_n254# 0.04fF
C11 a_1403_n44# w_n1957_n254# 0.04fF
C12 a_1045_n44# w_n1957_n254# 0.04fF
C13 a_687_n44# w_n1957_n254# 0.04fF
C14 a_329_n44# w_n1957_n254# 0.04fF
C15 a_n29_n44# w_n1957_n254# 0.04fF
C16 a_n387_n44# w_n1957_n254# 0.04fF
C17 a_n745_n44# w_n1957_n254# 0.04fF
C18 a_n1103_n44# w_n1957_n254# 0.04fF
C19 a_n1461_n44# w_n1957_n254# 0.04fF
C20 a_n1819_n44# w_n1957_n254# 0.04fF
C21 a_n1761_n132# w_n1957_n254# 3.23fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ND88ZC VSUBS a_303_n150# a_n753_n150# a_n369_n150#
+ w_n1367_n369# a_207_n150# a_n657_n150# a_591_n150# a_n1229_n150# a_n945_n150# a_495_n150#
+ a_n1041_n150# a_n849_n150# a_n81_n150# a_399_n150# a_783_n150# a_1071_n150# a_687_n150#
+ a_975_n150# a_n1137_n150# a_n273_n150# a_111_n150# a_879_n150# a_n177_n150# a_n561_n150#
+ a_15_n150# a_1167_n150# a_n1167_n247# a_n465_n150#
X0 a_n1137_n150# a_n1167_n247# a_n1229_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_495_n150# a_n1167_n247# a_399_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n561_n150# a_n1167_n247# a_n657_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_111_n150# a_n1167_n247# a_15_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_783_n150# a_n1167_n247# a_687_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_1071_n150# a_n1167_n247# a_975_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_399_n150# a_n1167_n247# a_303_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n465_n150# a_n1167_n247# a_n561_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_687_n150# a_n1167_n247# a_591_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n753_n150# a_n1167_n247# a_n849_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_975_n150# a_n1167_n247# a_879_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n81_n150# a_n1167_n247# a_n177_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_15_n150# a_n1167_n247# a_n81_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_n1041_n150# a_n1167_n247# a_n1137_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n369_n150# a_n1167_n247# a_n465_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_n657_n150# a_n1167_n247# a_n753_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_879_n150# a_n1167_n247# a_783_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_n945_n150# a_n1167_n247# a_n1041_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_1167_n150# a_n1167_n247# a_1071_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_303_n150# a_n1167_n247# a_207_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X20 a_n273_n150# a_n1167_n247# a_n369_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X21 a_591_n150# a_n1167_n247# a_495_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X22 a_n849_n150# a_n1167_n247# a_n945_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_207_n150# a_n1167_n247# a_111_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X24 a_n177_n150# a_n1167_n247# a_n273_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_399_n150# a_207_n150# 0.16fF
C1 a_n657_n150# a_n849_n150# 0.16fF
C2 a_1167_n150# w_n1367_n369# 0.14fF
C3 a_n369_n150# a_15_n150# 0.07fF
C4 a_n1137_n150# a_n849_n150# 0.10fF
C5 a_n177_n150# a_207_n150# 0.07fF
C6 a_111_n150# a_303_n150# 0.16fF
C7 a_495_n150# a_303_n150# 0.16fF
C8 a_111_n150# a_207_n150# 0.43fF
C9 a_399_n150# a_783_n150# 0.07fF
C10 a_n177_n150# a_n273_n150# 0.43fF
C11 a_495_n150# a_207_n150# 0.10fF
C12 a_n657_n150# a_n753_n150# 0.43fF
C13 a_687_n150# a_975_n150# 0.10fF
C14 a_111_n150# a_n273_n150# 0.07fF
C15 a_n1137_n150# a_n1229_n150# 0.43fF
C16 a_879_n150# a_783_n150# 0.43fF
C17 a_975_n150# a_591_n150# 0.07fF
C18 a_975_n150# w_n1367_n369# 0.05fF
C19 a_n1137_n150# a_n753_n150# 0.07fF
C20 a_n81_n150# a_n369_n150# 0.10fF
C21 a_n1229_n150# a_n849_n150# 0.07fF
C22 a_n81_n150# a_n465_n150# 0.07fF
C23 a_303_n150# a_15_n150# 0.10fF
C24 a_207_n150# a_15_n150# 0.16fF
C25 a_1071_n150# a_783_n150# 0.10fF
C26 a_n753_n150# a_n849_n150# 0.43fF
C27 a_n273_n150# a_15_n150# 0.10fF
C28 a_495_n150# a_783_n150# 0.10fF
C29 a_111_n150# a_399_n150# 0.10fF
C30 a_879_n150# a_1071_n150# 0.16fF
C31 a_495_n150# a_399_n150# 0.43fF
C32 a_n1041_n150# a_n945_n150# 0.43fF
C33 a_1167_n150# a_783_n150# 0.07fF
C34 a_n81_n150# a_303_n150# 0.07fF
C35 a_687_n150# a_591_n150# 0.43fF
C36 a_495_n150# a_879_n150# 0.07fF
C37 a_n81_n150# a_207_n150# 0.10fF
C38 a_n561_n150# a_n945_n150# 0.07fF
C39 a_n81_n150# a_n273_n150# 0.16fF
C40 a_879_n150# a_1167_n150# 0.10fF
C41 a_n177_n150# a_111_n150# 0.10fF
C42 a_399_n150# a_15_n150# 0.07fF
C43 a_n465_n150# a_n369_n150# 0.43fF
C44 a_n561_n150# a_n369_n150# 0.16fF
C45 a_495_n150# a_111_n150# 0.07fF
C46 a_n465_n150# a_n561_n150# 0.43fF
C47 a_975_n150# a_783_n150# 0.16fF
C48 a_1071_n150# a_1167_n150# 0.43fF
C49 a_687_n150# a_303_n150# 0.07fF
C50 a_n177_n150# a_15_n150# 0.16fF
C51 a_591_n150# a_303_n150# 0.10fF
C52 a_111_n150# a_15_n150# 0.43fF
C53 a_591_n150# a_207_n150# 0.07fF
C54 a_879_n150# a_975_n150# 0.43fF
C55 a_n657_n150# a_n945_n150# 0.10fF
C56 a_n273_n150# a_n369_n150# 0.43fF
C57 a_n1137_n150# a_n945_n150# 0.16fF
C58 a_n657_n150# a_n1041_n150# 0.07fF
C59 a_n465_n150# a_n273_n150# 0.16fF
C60 a_n657_n150# a_n369_n150# 0.10fF
C61 a_1071_n150# a_975_n150# 0.43fF
C62 a_n561_n150# a_n273_n150# 0.10fF
C63 a_n177_n150# a_n81_n150# 0.43fF
C64 a_n657_n150# a_n465_n150# 0.16fF
C65 a_n1137_n150# a_n1041_n150# 0.43fF
C66 a_n849_n150# a_n945_n150# 0.43fF
C67 a_687_n150# a_783_n150# 0.43fF
C68 a_n657_n150# a_n561_n150# 0.43fF
C69 a_111_n150# a_n81_n150# 0.16fF
C70 a_591_n150# a_783_n150# 0.16fF
C71 a_687_n150# a_399_n150# 0.10fF
C72 a_n1041_n150# a_n849_n150# 0.16fF
C73 a_303_n150# a_207_n150# 0.43fF
C74 a_399_n150# a_591_n150# 0.16fF
C75 a_879_n150# a_687_n150# 0.16fF
C76 a_975_n150# a_1167_n150# 0.16fF
C77 a_n1229_n150# a_n945_n150# 0.10fF
C78 a_n465_n150# a_n849_n150# 0.07fF
C79 a_879_n150# a_591_n150# 0.10fF
C80 a_n561_n150# a_n849_n150# 0.10fF
C81 a_879_n150# w_n1367_n369# 0.04fF
C82 a_n753_n150# a_n945_n150# 0.16fF
C83 a_n81_n150# a_15_n150# 0.43fF
C84 a_n1041_n150# a_n1229_n150# 0.16fF
C85 a_687_n150# a_1071_n150# 0.07fF
C86 a_n753_n150# a_n1041_n150# 0.10fF
C87 a_n657_n150# a_n273_n150# 0.07fF
C88 a_n753_n150# a_n369_n150# 0.07fF
C89 a_1071_n150# w_n1367_n369# 0.07fF
C90 a_495_n150# a_687_n150# 0.16fF
C91 a_n177_n150# a_n369_n150# 0.16fF
C92 a_n465_n150# a_n753_n150# 0.10fF
C93 a_n177_n150# a_n465_n150# 0.10fF
C94 a_495_n150# a_591_n150# 0.43fF
C95 a_n753_n150# a_n561_n150# 0.16fF
C96 a_399_n150# a_303_n150# 0.43fF
C97 a_n177_n150# a_n561_n150# 0.07fF
C98 a_1167_n150# VSUBS 0.03fF
C99 a_1071_n150# VSUBS 0.03fF
C100 a_975_n150# VSUBS 0.03fF
C101 a_879_n150# VSUBS 0.03fF
C102 a_783_n150# VSUBS 0.03fF
C103 a_687_n150# VSUBS 0.03fF
C104 a_591_n150# VSUBS 0.03fF
C105 a_495_n150# VSUBS 0.03fF
C106 a_399_n150# VSUBS 0.03fF
C107 a_303_n150# VSUBS 0.03fF
C108 a_207_n150# VSUBS 0.03fF
C109 a_111_n150# VSUBS 0.03fF
C110 a_15_n150# VSUBS 0.03fF
C111 a_n81_n150# VSUBS 0.03fF
C112 a_n177_n150# VSUBS 0.03fF
C113 a_n273_n150# VSUBS 0.03fF
C114 a_n369_n150# VSUBS 0.03fF
C115 a_n465_n150# VSUBS 0.03fF
C116 a_n561_n150# VSUBS 0.03fF
C117 a_n657_n150# VSUBS 0.03fF
C118 a_n753_n150# VSUBS 0.03fF
C119 a_n849_n150# VSUBS 0.03fF
C120 a_n945_n150# VSUBS 0.03fF
C121 a_n1041_n150# VSUBS 0.03fF
C122 a_n1137_n150# VSUBS 0.03fF
C123 a_n1229_n150# VSUBS 0.03fF
C124 a_n1167_n247# VSUBS 2.63fF
C125 w_n1367_n369# VSUBS 7.85fF
.ends

.subckt charge_pump vss pswitch nswitch out vdd biasp nUp Down w_2544_775# iref nDown
+ Up w_1008_774#
Xsky130_fd_pr__pfet_01v8_4ML9WA_0 vss pswitch vdd pswitch pswitch pswitch nUp pswitch
+ pswitch pswitch pswitch pswitch pswitch pswitch sky130_fd_pr__pfet_01v8_4ML9WA
Xsky130_fd_pr__nfet_01v8_YCGG98_0 vss out out vss vss vss out out vss vss out vss
+ out out out vss out vss out out out vss vss vss out vss vss nswitch sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_1 iref vss vss iref iref iref vss vss iref iref vss
+ iref vss vss vss iref vss iref vss vss vss vss iref iref vss iref iref iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_2 biasp vss vss biasp biasp biasp vss vss biasp biasp
+ vss biasp vss vss vss biasp vss biasp vss vss vss vss biasp biasp vss biasp biasp
+ iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_MUHGM9_0 nDown iref nswitch vss nswitch nswitch vss nswitch
+ iref nswitch nswitch vss nswitch Down iref iref vss vss nswitch nswitch iref nswitch
+ vss nswitch sky130_fd_pr__nfet_01v8_MUHGM9
Xsky130_fd_pr__pfet_01v8_NKZXKB_0 vss Up pswitch pswitch pswitch vdd biasp pswitch
+ pswitch pswitch vdd vdd biasp pswitch pswitch nUp vdd biasp pswitch pswitch vdd
+ pswitch biasp biasp vdd sky130_fd_pr__pfet_01v8_NKZXKB
Xsky130_fd_pr__nfet_01v8_8GRULZ_0 Down nswitch nswitch nswitch nswitch nswitch nswitch
+ nswitch nswitch nswitch vss nswitch nswitch sky130_fd_pr__nfet_01v8_8GRULZ
Xsky130_fd_pr__pfet_01v8_ND88ZC_0 vss vdd out out vdd out vdd out vdd out vdd vdd
+ vdd vdd out out vdd vdd out out vdd vdd vdd out out out out pswitch vdd sky130_fd_pr__pfet_01v8_ND88ZC
Xsky130_fd_pr__pfet_01v8_ND88ZC_1 vss biasp vdd vdd vdd vdd biasp vdd biasp vdd biasp
+ biasp biasp biasp vdd vdd biasp biasp vdd vdd biasp biasp biasp vdd vdd vdd vdd
+ biasp biasp sky130_fd_pr__pfet_01v8_ND88ZC
C0 Down nswitch 2.27fF
C1 Up nUp 0.15fF
C2 pswitch Up 0.70fF
C3 pswitch nUp 5.66fF
C4 pswitch biasp 3.11fF
C5 Down nUp 0.25fF
C6 out vdd 6.66fF
C7 nDown nswitch 0.31fF
C8 iref nswitch 1.91fF
C9 nswitch vdd 0.07fF
C10 out nswitch 1.28fF
C11 iref biasp 0.80fF
C12 vdd biasp 2.64fF
C13 out nUp 0.31fF
C14 pswitch vdd 3.98fF
C15 nDown Down 0.13fF
C16 pswitch out 4.91fF
C17 nswitch biasp 0.03fF
C18 pswitch nswitch 0.06fF
C19 vdd vss 35.71fF
C20 Down vss 4.77fF
C21 Up vss 1.17fF
C22 nswitch vss 6.39fF
C23 nDown vss 1.11fF
C24 biasp vss 8.73fF
C25 iref vss 10.12fF
C26 out vss -3.49fF
C27 pswitch vss 3.45fF
C28 nUp vss 5.85fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4798MH VSUBS a_81_n156# a_111_n125# a_15_n125# a_n173_n125#
+ w_n311_n344# a_n111_n156# a_n15_n156# a_n81_n125#
X0 a_n81_n125# a_n111_n156# a_n173_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n15_n156# a_n81_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_81_n156# a_15_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 w_n311_n344# a_n81_n125# 0.09fF
C1 a_n173_n125# a_n81_n125# 0.36fF
C2 a_111_n125# w_n311_n344# 0.14fF
C3 a_111_n125# a_n173_n125# 0.08fF
C4 a_111_n125# a_n81_n125# 0.13fF
C5 a_81_n156# a_n15_n156# 0.02fF
C6 w_n311_n344# a_15_n125# 0.09fF
C7 a_15_n125# a_n173_n125# 0.13fF
C8 w_n311_n344# a_n173_n125# 0.14fF
C9 a_15_n125# a_n81_n125# 0.36fF
C10 a_n111_n156# a_n15_n156# 0.02fF
C11 a_111_n125# a_15_n125# 0.36fF
C12 a_111_n125# VSUBS 0.03fF
C13 a_15_n125# VSUBS 0.03fF
C14 a_n81_n125# VSUBS 0.03fF
C15 a_n173_n125# VSUBS 0.03fF
C16 a_81_n156# VSUBS 0.05fF
C17 a_n15_n156# VSUBS 0.05fF
C18 a_n111_n156# VSUBS 0.05fF
C19 w_n311_n344# VSUBS 2.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_BHR94T a_n15_n151# w_n311_n335# a_81_n151# a_111_n125#
+ a_15_n125# a_n173_n125# a_n111_n151# a_n81_n125#
X0 a_111_n125# a_81_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n15_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_15_n125# a_n81_n125# 0.36fF
C1 a_15_n125# a_111_n125# 0.36fF
C2 a_n173_n125# a_n81_n125# 0.36fF
C3 a_n15_n151# a_81_n151# 0.02fF
C4 a_n173_n125# a_111_n125# 0.08fF
C5 a_n15_n151# a_n111_n151# 0.02fF
C6 a_n173_n125# a_15_n125# 0.13fF
C7 a_111_n125# a_n81_n125# 0.13fF
C8 a_111_n125# w_n311_n335# 0.17fF
C9 a_15_n125# w_n311_n335# 0.12fF
C10 a_n81_n125# w_n311_n335# 0.12fF
C11 a_n173_n125# w_n311_n335# 0.17fF
C12 a_81_n151# w_n311_n335# 0.05fF
C13 a_n15_n151# w_n311_n335# 0.05fF
C14 a_n111_n151# w_n311_n335# 0.05fF
.ends

.subckt trans_gate m1_187_n605# m1_45_n513# vss vdd
Xsky130_fd_pr__pfet_01v8_4798MH_0 vss vss m1_187_n605# m1_45_n513# m1_45_n513# vdd
+ vss vss m1_187_n605# sky130_fd_pr__pfet_01v8_4798MH
Xsky130_fd_pr__nfet_01v8_BHR94T_0 vdd vss vdd m1_187_n605# m1_45_n513# m1_45_n513#
+ vdd m1_187_n605# sky130_fd_pr__nfet_01v8_BHR94T
C0 m1_45_n513# m1_187_n605# 0.36fF
C1 m1_45_n513# vdd 0.69fF
C2 vdd m1_187_n605# 0.55fF
C3 m1_187_n605# vss 0.93fF
C4 m1_45_n513# vss 1.31fF
C5 vdd vss 3.36fF
.ends

.subckt sky130_fd_pr__pfet_01v8_7KT7MH VSUBS a_n111_n186# a_111_n125# a_15_n125# a_n173_n125#
+ w_n311_n344# a_n81_n125#
X0 a_n81_n125# a_n111_n186# a_n173_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n111_n186# a_n81_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_n111_n186# a_15_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_111_n125# w_n311_n344# 0.14fF
C1 a_n173_n125# a_n81_n125# 0.36fF
C2 a_n173_n125# a_15_n125# 0.13fF
C3 a_111_n125# a_n173_n125# 0.08fF
C4 a_15_n125# a_n81_n125# 0.36fF
C5 a_n173_n125# w_n311_n344# 0.14fF
C6 a_111_n125# a_n81_n125# 0.13fF
C7 a_n81_n125# w_n311_n344# 0.09fF
C8 a_111_n125# a_15_n125# 0.36fF
C9 a_15_n125# w_n311_n344# 0.09fF
C10 a_111_n125# VSUBS 0.03fF
C11 a_15_n125# VSUBS 0.03fF
C12 a_n81_n125# VSUBS 0.03fF
C13 a_n173_n125# VSUBS 0.03fF
C14 a_n111_n186# VSUBS 0.26fF
C15 w_n311_n344# VSUBS 2.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS6QM w_n311_n335# a_111_n125# a_15_n125# a_n173_n125#
+ a_n111_n151# a_n81_n125#
X0 a_111_n125# a_n111_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n111_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n81_n125# a_15_n125# 0.36fF
C1 a_n81_n125# a_111_n125# 0.13fF
C2 a_n173_n125# a_n81_n125# 0.36fF
C3 a_111_n125# a_15_n125# 0.36fF
C4 a_n173_n125# a_15_n125# 0.13fF
C5 a_n173_n125# a_111_n125# 0.08fF
C6 a_111_n125# w_n311_n335# 0.17fF
C7 a_15_n125# w_n311_n335# 0.12fF
C8 a_n81_n125# w_n311_n335# 0.12fF
C9 a_n173_n125# w_n311_n335# 0.17fF
C10 a_n111_n151# w_n311_n335# 0.25fF
.ends

.subckt inverter_cp_x1 out in vss vdd
Xsky130_fd_pr__pfet_01v8_7KT7MH_0 vss in out vdd vdd vdd out sky130_fd_pr__pfet_01v8_7KT7MH
Xsky130_fd_pr__nfet_01v8_2BS6QM_0 vss out vss vss in out sky130_fd_pr__nfet_01v8_2BS6QM
C0 out vdd 0.10fF
C1 out in 0.32fF
C2 out vss 0.77fF
C3 in vss 0.95fF
C4 vdd vss 3.13fF
.ends

.subckt clock_inverter vss inverter_cp_x1_2/in CLK vdd inverter_cp_x1_0/out CLK_d
+ nCLK_d
Xtrans_gate_0 nCLK_d inverter_cp_x1_0/out vss vdd trans_gate
Xinverter_cp_x1_0 inverter_cp_x1_0/out CLK vss vdd inverter_cp_x1
Xinverter_cp_x1_1 inverter_cp_x1_2/in CLK vss vdd inverter_cp_x1
Xinverter_cp_x1_2 CLK_d inverter_cp_x1_2/in vss vdd inverter_cp_x1
C0 nCLK_d vdd 0.03fF
C1 inverter_cp_x1_2/in vdd 0.21fF
C2 inverter_cp_x1_0/out CLK 0.31fF
C3 inverter_cp_x1_0/out nCLK_d 0.11fF
C4 inverter_cp_x1_2/in CLK_d 0.12fF
C5 inverter_cp_x1_2/in CLK 0.31fF
C6 inverter_cp_x1_0/out vdd 0.28fF
C7 CLK_d vdd 0.03fF
C8 CLK vdd 0.36fF
C9 CLK_d vss 0.96fF
C10 inverter_cp_x1_2/in vss 2.01fF
C11 inverter_cp_x1_0/out vss 1.97fF
C12 CLK vss 3.03fF
C13 nCLK_d vss 1.44fF
C14 vdd vss 16.51fF
.ends

.subckt sky130_fd_pr__pfet_01v8_MJG8BZ VSUBS a_n125_n95# a_63_n95# w_n263_n314# a_n33_n95#
+ a_n63_n192#
X0 a_63_n95# a_n63_n192# a_n33_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n33_n95# a_n63_n192# a_n125_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
C0 a_n125_n95# a_n33_n95# 0.28fF
C1 a_n125_n95# w_n263_n314# 0.11fF
C2 w_n263_n314# a_n33_n95# 0.08fF
C3 a_n125_n95# a_63_n95# 0.10fF
C4 a_63_n95# a_n33_n95# 0.28fF
C5 a_63_n95# w_n263_n314# 0.11fF
C6 a_63_n95# VSUBS 0.03fF
C7 a_n33_n95# VSUBS 0.03fF
C8 a_n125_n95# VSUBS 0.03fF
C9 a_n63_n192# VSUBS 0.20fF
C10 w_n263_n314# VSUBS 1.80fF
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS854 w_n311_n335# a_n129_n213# a_111_n125# a_15_n125#
+ a_n173_n125# a_n81_n125#
X0 a_111_n125# a_n129_n213# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n129_n213# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n129_n213# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_n173_n125# a_n129_n213# 0.02fF
C1 a_n81_n125# a_15_n125# 0.36fF
C2 a_n81_n125# a_n129_n213# 0.10fF
C3 a_n129_n213# a_15_n125# 0.10fF
C4 a_n173_n125# a_111_n125# 0.08fF
C5 a_n81_n125# a_111_n125# 0.13fF
C6 a_n173_n125# a_n81_n125# 0.36fF
C7 a_111_n125# a_15_n125# 0.36fF
C8 a_111_n125# a_n129_n213# 0.01fF
C9 a_n173_n125# a_15_n125# 0.13fF
C10 a_111_n125# w_n311_n335# 0.05fF
C11 a_15_n125# w_n311_n335# 0.05fF
C12 a_n81_n125# w_n311_n335# 0.05fF
C13 a_n173_n125# w_n311_n335# 0.05fF
C14 a_n129_n213# w_n311_n335# 0.49fF
.ends

.subckt sky130_fd_pr__nfet_01v8_KU9PSX a_n125_n95# a_n33_n95# a_n81_n183# w_n263_n305#
X0 a_n33_n95# a_n81_n183# a_n125_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n125_n95# a_n81_n183# a_n33_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
C0 a_n125_n95# a_n81_n183# 0.16fF
C1 a_n33_n95# a_n81_n183# 0.10fF
C2 a_n125_n95# a_n33_n95# 0.88fF
C3 a_n33_n95# w_n263_n305# 0.07fF
C4 a_n125_n95# w_n263_n305# 0.13fF
C5 a_n81_n183# w_n263_n305# 0.31fF
.ends

.subckt latch_diff m1_657_280# nQ Q vss CLK vdd nD D
Xsky130_fd_pr__pfet_01v8_MJG8BZ_0 vss vdd vdd vdd nQ Q sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__pfet_01v8_MJG8BZ_1 vss vdd vdd vdd Q nQ sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__nfet_01v8_2BS854_0 vss CLK vss m1_657_280# m1_657_280# vss sky130_fd_pr__nfet_01v8_2BS854
Xsky130_fd_pr__nfet_01v8_KU9PSX_0 m1_657_280# Q nD vss sky130_fd_pr__nfet_01v8_KU9PSX
Xsky130_fd_pr__nfet_01v8_KU9PSX_1 m1_657_280# nQ D vss sky130_fd_pr__nfet_01v8_KU9PSX
C0 m1_657_280# CLK 0.24fF
C1 m1_657_280# Q 0.94fF
C2 nQ D 0.05fF
C3 nQ m1_657_280# 1.41fF
C4 nD Q 0.05fF
C5 nQ Q 0.93fF
C6 vdd Q 0.16fF
C7 nQ nD 0.05fF
C8 Q D 0.05fF
C9 nQ vdd 0.16fF
C10 nQ vss 1.16fF
C11 D vss 0.53fF
C12 Q vss -0.55fF
C13 m1_657_280# vss 1.88fF
C14 nD vss 0.16fF
C15 CLK vss 0.87fF
C16 vdd vss 5.98fF
.ends

.subckt DFlipFlop latch_diff_0/m1_657_280# vss latch_diff_1/D clock_inverter_0/inverter_cp_x1_2/in
+ nQ Q latch_diff_1/nD D latch_diff_1/m1_657_280# latch_diff_0/D vdd CLK clock_inverter_0/inverter_cp_x1_0/out
+ nCLK latch_diff_0/nD
Xclock_inverter_0 vss clock_inverter_0/inverter_cp_x1_2/in D vdd clock_inverter_0/inverter_cp_x1_0/out
+ latch_diff_0/D latch_diff_0/nD clock_inverter
Xlatch_diff_0 latch_diff_0/m1_657_280# latch_diff_1/nD latch_diff_1/D vss CLK vdd
+ latch_diff_0/nD latch_diff_0/D latch_diff
Xlatch_diff_1 latch_diff_1/m1_657_280# nQ Q vss nCLK vdd latch_diff_1/nD latch_diff_1/D
+ latch_diff
C0 latch_diff_1/D latch_diff_1/m1_657_280# 0.32fF
C1 clock_inverter_0/inverter_cp_x1_0/out vdd 0.03fF
C2 latch_diff_1/D latch_diff_0/nD 0.41fF
C3 latch_diff_1/D nQ 0.11fF
C4 latch_diff_1/nD latch_diff_0/m1_657_280# 0.14fF
C5 latch_diff_0/D latch_diff_0/m1_657_280# 0.37fF
C6 latch_diff_1/nD vdd 0.02fF
C7 latch_diff_1/nD latch_diff_0/D 0.04fF
C8 latch_diff_1/m1_657_280# latch_diff_0/m1_657_280# 0.18fF
C9 vdd latch_diff_0/D 0.09fF
C10 latch_diff_1/nD latch_diff_1/m1_657_280# 0.42fF
C11 latch_diff_0/m1_657_280# latch_diff_0/nD 0.38fF
C12 Q latch_diff_1/nD 0.01fF
C13 nQ latch_diff_1/nD 0.08fF
C14 latch_diff_1/D latch_diff_0/m1_657_280# 0.43fF
C15 vdd latch_diff_0/nD 0.14fF
C16 latch_diff_1/D latch_diff_1/nD 0.33fF
C17 latch_diff_1/D vdd 0.03fF
C18 latch_diff_1/D latch_diff_0/D 0.11fF
C19 nQ vss 0.57fF
C20 Q vss -0.92fF
C21 latch_diff_1/m1_657_280# vss 0.64fF
C22 nCLK vss 0.83fF
C23 latch_diff_1/nD vss 1.83fF
C24 latch_diff_1/D vss -0.30fF
C25 latch_diff_0/m1_657_280# vss 0.72fF
C26 CLK vss 0.83fF
C27 latch_diff_0/D vss 1.29fF
C28 clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C29 clock_inverter_0/inverter_cp_x1_0/out vss 1.84fF
C30 D vss 3.27fF
C31 latch_diff_0/nD vss 1.74fF
C32 vdd vss 32.62fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ZP3U9B VSUBS a_n221_n84# a_159_n84# w_n359_n303# a_n63_n110#
+ a_n129_n84# a_33_n110# a_n159_n110# a_63_n84# a_129_n110# a_n33_n84#
X0 a_n129_n84# a_n159_n110# a_n221_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_63_n84# a_33_n110# a_n33_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_n33_n84# a_n63_n110# a_n129_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_159_n84# a_129_n110# a_63_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_33_n110# a_129_n110# 0.02fF
C1 a_n221_n84# a_159_n84# 0.04fF
C2 a_n221_n84# a_n33_n84# 0.09fF
C3 a_n63_n110# a_n159_n110# 0.02fF
C4 a_n221_n84# a_n129_n84# 0.24fF
C5 w_n359_n303# a_n221_n84# 0.08fF
C6 a_n33_n84# a_159_n84# 0.09fF
C7 a_n129_n84# a_159_n84# 0.05fF
C8 w_n359_n303# a_159_n84# 0.08fF
C9 a_n33_n84# a_n129_n84# 0.24fF
C10 w_n359_n303# a_n33_n84# 0.05fF
C11 w_n359_n303# a_n129_n84# 0.06fF
C12 a_n221_n84# a_63_n84# 0.05fF
C13 a_63_n84# a_159_n84# 0.24fF
C14 a_n63_n110# a_33_n110# 0.02fF
C15 a_n33_n84# a_63_n84# 0.24fF
C16 a_63_n84# a_n129_n84# 0.09fF
C17 w_n359_n303# a_63_n84# 0.06fF
C18 a_159_n84# VSUBS 0.03fF
C19 a_63_n84# VSUBS 0.03fF
C20 a_n33_n84# VSUBS 0.03fF
C21 a_n129_n84# VSUBS 0.03fF
C22 a_n221_n84# VSUBS 0.03fF
C23 a_129_n110# VSUBS 0.05fF
C24 a_33_n110# VSUBS 0.05fF
C25 a_n63_n110# VSUBS 0.05fF
C26 a_n159_n110# VSUBS 0.05fF
C27 w_n359_n303# VSUBS 2.19fF
.ends

.subckt sky130_fd_pr__nfet_01v8_DXA56D w_n359_n252# a_n33_n42# a_129_n68# a_n159_n68#
+ a_n221_n42# a_159_n42# a_n129_n42# a_33_n68# a_n63_n68# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n129_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_159_n42# a_129_n68# a_63_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_n129_n42# a_n159_n68# a_n221_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n221_n42# a_n33_n42# 0.05fF
C1 a_159_n42# a_63_n42# 0.12fF
C2 a_159_n42# a_n221_n42# 0.02fF
C3 a_63_n42# a_n129_n42# 0.05fF
C4 a_159_n42# a_n33_n42# 0.05fF
C5 a_n221_n42# a_n129_n42# 0.12fF
C6 a_33_n68# a_n63_n68# 0.02fF
C7 a_n33_n42# a_n129_n42# 0.12fF
C8 a_n159_n68# a_n63_n68# 0.02fF
C9 a_n221_n42# a_63_n42# 0.03fF
C10 a_129_n68# a_33_n68# 0.02fF
C11 a_63_n42# a_n33_n42# 0.12fF
C12 a_159_n42# a_n129_n42# 0.03fF
C13 a_159_n42# w_n359_n252# 0.07fF
C14 a_63_n42# w_n359_n252# 0.06fF
C15 a_n33_n42# w_n359_n252# 0.06fF
C16 a_n129_n42# w_n359_n252# 0.06fF
C17 a_n221_n42# w_n359_n252# 0.07fF
C18 a_129_n68# w_n359_n252# 0.05fF
C19 a_33_n68# w_n359_n252# 0.05fF
C20 a_n63_n68# w_n359_n252# 0.05fF
C21 a_n159_n68# w_n359_n252# 0.05fF
.ends

.subckt inverter_min_x4 in vss out vdd
Xsky130_fd_pr__pfet_01v8_ZP3U9B_0 vss out out vdd in vdd in in vdd in out sky130_fd_pr__pfet_01v8_ZP3U9B
Xsky130_fd_pr__nfet_01v8_DXA56D_0 vss out in in out out vss in in vss sky130_fd_pr__nfet_01v8_DXA56D
C0 vdd out 0.62fF
C1 in out 0.67fF
C2 in vdd 0.33fF
C3 out vss 0.66fF
C4 in vss 1.89fF
C5 vdd vss 3.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_5RJ8EK a_n33_n42# a_33_n68# w_n263_n252# a_n63_n68#
+ a_n125_n42# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n125_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n33_n42# a_n125_n42# 0.12fF
C1 a_n63_n68# a_33_n68# 0.02fF
C2 a_n125_n42# a_63_n42# 0.05fF
C3 a_n33_n42# a_63_n42# 0.12fF
C4 a_63_n42# w_n263_n252# 0.09fF
C5 a_n33_n42# w_n263_n252# 0.07fF
C6 a_n125_n42# w_n263_n252# 0.09fF
C7 a_33_n68# w_n263_n252# 0.05fF
C8 a_n63_n68# w_n263_n252# 0.05fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ZPB9BB VSUBS a_n63_n110# a_33_n110# a_n125_n84# a_63_n84#
+ w_n263_n303# a_n33_n84#
X0 a_63_n84# a_33_n110# a_n33_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_n33_n84# a_n63_n110# a_n125_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_n125_n84# a_63_n84# 0.09fF
C1 a_n125_n84# w_n263_n303# 0.10fF
C2 a_33_n110# a_n63_n110# 0.02fF
C3 a_63_n84# a_n33_n84# 0.24fF
C4 w_n263_n303# a_n33_n84# 0.07fF
C5 a_63_n84# w_n263_n303# 0.10fF
C6 a_n125_n84# a_n33_n84# 0.24fF
C7 a_63_n84# VSUBS 0.03fF
C8 a_n33_n84# VSUBS 0.03fF
C9 a_n125_n84# VSUBS 0.03fF
C10 a_33_n110# VSUBS 0.05fF
C11 a_n63_n110# VSUBS 0.05fF
C12 w_n263_n303# VSUBS 1.74fF
.ends

.subckt inverter_min_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_5RJ8EK_0 vss in vss in out out sky130_fd_pr__nfet_01v8_5RJ8EK
Xsky130_fd_pr__pfet_01v8_ZPB9BB_0 vss in in out out vdd vdd sky130_fd_pr__pfet_01v8_ZPB9BB
C0 vdd out 0.15fF
C1 vdd in 0.01fF
C2 out in 0.30fF
C3 vdd vss 2.93fF
C4 out vss 0.66fF
C5 in vss 0.72fF
.ends

.subckt div_by_2 vss vdd clock_inverter_0/inverter_cp_x1_2/in CLK_2 nCLK_2 o1 CLK
+ out_div o2 clock_inverter_0/inverter_cp_x1_0/out nout_div
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vss DFlipFlop_0/latch_diff_1/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ nout_div out_div DFlipFlop_0/latch_diff_1/nD nout_div DFlipFlop_0/latch_diff_1/m1_657_280#
+ DFlipFlop_0/latch_diff_0/D vdd DFlipFlop_0/CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_0/nCLK DFlipFlop_0/latch_diff_0/nD DFlipFlop
Xclock_inverter_0 vss clock_inverter_0/inverter_cp_x1_2/in CLK vdd clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_0/CLK DFlipFlop_0/nCLK clock_inverter
Xinverter_min_x4_0 o1 vss CLK_2 vdd inverter_min_x4
Xinverter_min_x4_1 o2 vss nCLK_2 vdd inverter_min_x4
Xinverter_min_x2_0 nout_div o2 vss vdd inverter_min_x2
Xinverter_min_x2_1 out_div o1 vss vdd inverter_min_x2
C0 nout_div out_div 0.22fF
C1 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vdd 0.03fF
C2 o2 nCLK_2 0.11fF
C3 DFlipFlop_0/latch_diff_1/m1_657_280# DFlipFlop_0/nCLK 0.26fF
C4 nout_div DFlipFlop_0/latch_diff_0/D 0.09fF
C5 DFlipFlop_0/latch_diff_0/m1_657_280# DFlipFlop_0/CLK 0.26fF
C6 DFlipFlop_0/latch_diff_0/nD DFlipFlop_0/CLK 0.12fF
C7 vdd out_div 0.03fF
C8 clock_inverter_0/inverter_cp_x1_0/out vdd 0.10fF
C9 o2 vdd 0.14fF
C10 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vdd 0.03fF
C11 DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/nCLK -0.09fF
C12 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_0/nCLK 0.46fF
C13 o1 vdd 0.14fF
C14 DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/CLK 0.11fF
C15 DFlipFlop_0/latch_diff_0/D DFlipFlop_0/nCLK 0.13fF
C16 nout_div vdd 0.16fF
C17 DFlipFlop_0/latch_diff_1/D nout_div 0.64fF
C18 o2 DFlipFlop_0/latch_diff_1/m1_657_280# 0.02fF
C19 nCLK_2 vdd 0.08fF
C20 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop_0/CLK 0.29fF
C21 o1 CLK_2 0.11fF
C22 o1 DFlipFlop_0/latch_diff_1/m1_657_280# 0.02fF
C23 nout_div DFlipFlop_0/nCLK 0.43fF
C24 nout_div DFlipFlop_0/latch_diff_0/nD 0.07fF
C25 DFlipFlop_0/latch_diff_0/m1_657_280# nout_div 0.24fF
C26 nout_div DFlipFlop_0/CLK 0.42fF
C27 DFlipFlop_0/nCLK vdd 0.30fF
C28 nout_div DFlipFlop_0/latch_diff_1/m1_657_280# 0.21fF
C29 DFlipFlop_0/latch_diff_1/D DFlipFlop_0/nCLK 0.08fF
C30 o1 out_div 0.01fF
C31 CLK_2 vdd 0.08fF
C32 nout_div DFlipFlop_0/latch_diff_1/nD 1.18fF
C33 DFlipFlop_0/CLK vdd 0.40fF
C34 DFlipFlop_0/latch_diff_1/D DFlipFlop_0/CLK -0.48fF
C35 nCLK_2 vss 1.08fF
C36 o2 vss 2.21fF
C37 CLK_2 vss 1.08fF
C38 o1 vss 2.21fF
C39 DFlipFlop_0/CLK vss 1.03fF
C40 clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C41 clock_inverter_0/inverter_cp_x1_0/out vss 1.85fF
C42 CLK vss 3.27fF
C43 DFlipFlop_0/nCLK vss 1.76fF
C44 out_div vss -0.77fF
C45 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.63fF
C46 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C47 DFlipFlop_0/latch_diff_1/D vss -1.72fF
C48 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C49 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C50 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.89fF
C51 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.80fF
C52 nout_div vss 4.41fF
C53 DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C54 vdd vss 64.43fF
.ends

.subckt sky130_fd_pr__pfet_01v8_58ZKDE VSUBS a_n257_n777# a_n129_n600# a_n221_n600#
+ w_n257_n702#
X0 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X1 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X2 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X3 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
C0 a_n129_n600# a_n221_n600# 7.87fF
C1 a_n129_n600# a_n257_n777# 0.29fF
C2 a_n257_n777# a_n221_n600# 0.25fF
C3 a_n129_n600# VSUBS 0.10fF
C4 a_n221_n600# VSUBS 0.25fF
C5 a_n257_n777# VSUBS 1.05fF
C6 w_n257_n702# VSUBS 2.16fF
.ends

.subckt sky130_fd_pr__nfet_01v8_T69Y3A a_n129_n300# a_n221_n300# w_n257_n327# a_n257_n404#
X0 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
C0 a_n257_n404# a_n129_n300# 0.30fF
C1 a_n257_n404# a_n221_n300# 0.21fF
C2 a_n221_n300# a_n129_n300# 4.05fF
C3 a_n129_n300# w_n257_n327# 0.11fF
C4 a_n221_n300# w_n257_n327# 0.25fF
C5 a_n257_n404# w_n257_n327# 1.11fF
.ends

.subckt buffer_salida a_678_n100# out in a_3996_n100# vss vdd
Xsky130_fd_pr__pfet_01v8_58ZKDE_1 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_2 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_3 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_0 a_678_n100# vss vss in sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_1 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_4 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_5 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_2 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_3 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_6 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_70 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_4 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_7 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_8 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_71 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_60 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_5 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_72 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_61 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_50 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_6 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_9 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_62 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_51 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_7 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_40 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_8 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_63 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_52 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_30 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_41 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_64 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_53 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_9 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_20 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_31 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_42 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_65 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_54 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_10 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_21 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_32 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_43 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_66 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_55 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_11 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_22 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_33 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_44 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_67 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_56 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_12 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_23 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_34 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_45 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_68 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_57 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_13 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_24 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_35 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_46 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_69 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_58 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_14 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_25 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_36 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_47 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_59 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_48 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_15 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_26 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_37 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_49 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_16 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_27 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_38 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_70 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_17 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_28 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_39 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_71 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_60 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_18 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_29 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_72 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_61 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_50 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_62 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_51 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_19 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_40 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_63 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_52 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_30 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_41 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_64 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_53 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_20 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_31 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_42 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_65 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_54 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_10 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_21 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_32 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_43 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_66 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_55 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_11 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_22 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_33 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_44 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_67 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_56 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_12 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_23 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_34 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_45 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_68 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_57 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_46 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_13 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_24 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_35 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_69 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_58 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_14 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_25 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_36 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_47 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_59 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_15 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_26 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_37 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_48 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_49 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_16 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_27 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_38 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_17 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_28 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_39 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_18 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_29 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_19 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_0 vss in a_678_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
C0 a_678_n100# vdd 0.08fF
C1 in vdd 0.02fF
C2 out vdd 47.17fF
C3 in a_678_n100# 0.81fF
C4 a_3996_n100# vdd 3.68fF
C5 a_3996_n100# a_678_n100# 6.52fF
C6 a_3996_n100# out 55.19fF
C7 vdd vss 20.93fF
C8 out vss 35.17fF
C9 a_3996_n100# vss 49.53fF
C10 a_678_n100# vss 13.08fF
C11 in vss 0.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_CBAU6Y a_n73_n150# a_n33_n238# w_n211_n360# a_15_n150#
X0 a_15_n150# a_n33_n238# a_n73_n150# w_n211_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n33_n238# a_15_n150# 0.02fF
C1 a_n73_n150# a_15_n150# 0.51fF
C2 a_n33_n238# a_n73_n150# 0.02fF
C3 a_15_n150# w_n211_n360# 0.23fF
C4 a_n73_n150# w_n211_n360# 0.23fF
C5 a_n33_n238# w_n211_n360# 0.17fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4757AC VSUBS a_n73_n150# a_n33_181# w_n211_n369# a_15_n150#
X0 a_15_n150# a_n33_181# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 w_n211_n369# a_n73_n150# 0.20fF
C1 a_n33_181# a_n73_n150# 0.01fF
C2 a_15_n150# w_n211_n369# 0.20fF
C3 a_15_n150# a_n33_181# 0.01fF
C4 w_n211_n369# a_n33_181# 0.05fF
C5 a_15_n150# a_n73_n150# 0.51fF
C6 a_15_n150# VSUBS 0.03fF
C7 a_n73_n150# VSUBS 0.03fF
C8 a_n33_181# VSUBS 0.13fF
C9 w_n211_n369# VSUBS 1.98fF
.ends

.subckt sky130_fd_pr__nfet_01v8_7H8F5S a_n465_172# a_n417_n150# a_351_n150# a_255_n150#
+ w_n647_n360# a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150#
X0 a_159_n150# a_n465_172# a_63_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n225_n150# a_n465_172# a_n321_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_447_n150# a_n465_172# a_351_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_63_n150# a_n465_172# a_n33_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n465_172# a_n225_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n465_172# a_n509_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n33_n150# a_n465_172# a_n129_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_351_n150# a_n465_172# a_255_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_255_n150# a_n465_172# a_159_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n321_n150# a_n465_172# a_n417_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_63_n150# a_159_n150# 0.43fF
C1 a_n465_172# a_n417_n150# 0.10fF
C2 a_255_n150# a_63_n150# 0.16fF
C3 a_n321_n150# a_63_n150# 0.07fF
C4 a_n129_n150# a_63_n150# 0.16fF
C5 a_n33_n150# a_351_n150# 0.07fF
C6 a_n465_172# a_351_n150# 0.10fF
C7 a_n33_n150# a_63_n150# 0.43fF
C8 a_447_n150# a_159_n150# 0.10fF
C9 a_255_n150# a_447_n150# 0.16fF
C10 a_n465_172# a_63_n150# 0.10fF
C11 a_n225_n150# a_n509_n150# 0.10fF
C12 a_255_n150# a_159_n150# 0.43fF
C13 a_n129_n150# a_159_n150# 0.10fF
C14 a_n509_n150# a_n417_n150# 0.43fF
C15 a_255_n150# a_n129_n150# 0.07fF
C16 a_n321_n150# a_n129_n150# 0.16fF
C17 a_n465_172# a_447_n150# 0.01fF
C18 a_n33_n150# a_159_n150# 0.16fF
C19 a_255_n150# a_n33_n150# 0.10fF
C20 a_n321_n150# a_n33_n150# 0.10fF
C21 a_n465_172# a_159_n150# 0.10fF
C22 a_n33_n150# a_n129_n150# 0.43fF
C23 a_255_n150# a_n465_172# 0.10fF
C24 a_n321_n150# a_n465_172# 0.10fF
C25 a_n465_172# a_n129_n150# 0.10fF
C26 a_n465_172# a_n33_n150# 0.10fF
C27 a_n225_n150# a_n417_n150# 0.16fF
C28 a_n321_n150# a_n509_n150# 0.16fF
C29 a_n225_n150# a_63_n150# 0.10fF
C30 a_n129_n150# a_n509_n150# 0.07fF
C31 a_n465_172# a_n509_n150# 0.01fF
C32 a_351_n150# a_63_n150# 0.10fF
C33 a_n225_n150# a_159_n150# 0.07fF
C34 a_n321_n150# a_n225_n150# 0.43fF
C35 a_n225_n150# a_n129_n150# 0.43fF
C36 a_n321_n150# a_n417_n150# 0.43fF
C37 a_351_n150# a_447_n150# 0.43fF
C38 a_n129_n150# a_n417_n150# 0.10fF
C39 a_447_n150# a_63_n150# 0.07fF
C40 a_n33_n150# a_n225_n150# 0.16fF
C41 a_351_n150# a_159_n150# 0.16fF
C42 a_n465_172# a_n225_n150# 0.10fF
C43 a_n33_n150# a_n417_n150# 0.07fF
C44 a_255_n150# a_351_n150# 0.43fF
C45 a_447_n150# w_n647_n360# 0.17fF
C46 a_351_n150# w_n647_n360# 0.10fF
C47 a_255_n150# w_n647_n360# 0.08fF
C48 a_159_n150# w_n647_n360# 0.07fF
C49 a_63_n150# w_n647_n360# 0.04fF
C50 a_n33_n150# w_n647_n360# 0.04fF
C51 a_n129_n150# w_n647_n360# 0.04fF
C52 a_n225_n150# w_n647_n360# 0.07fF
C53 a_n321_n150# w_n647_n360# 0.08fF
C54 a_n417_n150# w_n647_n360# 0.10fF
C55 a_n509_n150# w_n647_n360# 0.17fF
C56 a_n465_172# w_n647_n360# 1.49fF
.ends

.subckt sky130_fd_pr__pfet_01v8_8DL6ZL VSUBS a_n417_n150# a_351_n150# a_255_n150#
+ a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n465_n247# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150# w_n647_n369#
X0 a_63_n150# a_n465_n247# a_n33_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n129_n150# a_n465_n247# a_n225_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n417_n150# a_n465_n247# a_n509_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n33_n150# a_n465_n247# a_n129_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_351_n150# a_n465_n247# a_255_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_255_n150# a_n465_n247# a_159_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n321_n150# a_n465_n247# a_n417_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_159_n150# a_n465_n247# a_63_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n225_n150# a_n465_n247# a_n321_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_447_n150# a_n465_n247# a_351_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
C0 a_n33_n150# a_63_n150# 0.43fF
C1 a_n33_n150# a_n129_n150# 0.43fF
C2 a_63_n150# a_n129_n150# 0.16fF
C3 a_n509_n150# a_n225_n150# 0.10fF
C4 a_n33_n150# a_159_n150# 0.16fF
C5 a_63_n150# a_159_n150# 0.43fF
C6 a_n321_n150# a_n417_n150# 0.43fF
C7 a_n33_n150# a_351_n150# 0.07fF
C8 a_159_n150# a_n129_n150# 0.10fF
C9 a_351_n150# a_63_n150# 0.10fF
C10 a_351_n150# a_159_n150# 0.16fF
C11 a_255_n150# a_447_n150# 0.16fF
C12 a_n321_n150# w_n647_n369# 0.05fF
C13 a_n417_n150# w_n647_n369# 0.07fF
C14 a_n465_n247# a_n321_n150# 0.08fF
C15 a_n465_n247# a_n417_n150# 0.08fF
C16 a_n321_n150# a_n225_n150# 0.43fF
C17 a_n225_n150# a_n417_n150# 0.16fF
C18 a_n465_n247# w_n647_n369# 0.47fF
C19 a_63_n150# a_447_n150# 0.07fF
C20 a_n225_n150# w_n647_n369# 0.04fF
C21 a_159_n150# a_447_n150# 0.10fF
C22 a_n465_n247# a_n225_n150# 0.08fF
C23 a_351_n150# a_447_n150# 0.43fF
C24 a_n509_n150# a_n129_n150# 0.07fF
C25 a_255_n150# w_n647_n369# 0.05fF
C26 a_n465_n247# a_255_n150# 0.08fF
C27 a_n33_n150# a_n321_n150# 0.10fF
C28 a_63_n150# a_n321_n150# 0.07fF
C29 a_n33_n150# a_n417_n150# 0.07fF
C30 a_n321_n150# a_n129_n150# 0.16fF
C31 a_n417_n150# a_n129_n150# 0.10fF
C32 a_n33_n150# w_n647_n369# 0.02fF
C33 a_63_n150# w_n647_n369# 0.02fF
C34 a_n129_n150# w_n647_n369# 0.02fF
C35 a_n465_n247# a_n33_n150# 0.08fF
C36 a_n465_n247# a_63_n150# 0.08fF
C37 a_n465_n247# a_n129_n150# 0.08fF
C38 a_159_n150# w_n647_n369# 0.04fF
C39 a_351_n150# w_n647_n369# 0.07fF
C40 a_n465_n247# a_159_n150# 0.08fF
C41 a_n33_n150# a_n225_n150# 0.16fF
C42 a_63_n150# a_n225_n150# 0.10fF
C43 a_n465_n247# a_351_n150# 0.08fF
C44 a_n225_n150# a_n129_n150# 0.43fF
C45 a_n225_n150# a_159_n150# 0.07fF
C46 a_447_n150# w_n647_n369# 0.14fF
C47 a_n33_n150# a_255_n150# 0.10fF
C48 a_63_n150# a_255_n150# 0.16fF
C49 a_255_n150# a_n129_n150# 0.07fF
C50 a_n509_n150# a_n321_n150# 0.16fF
C51 a_n509_n150# a_n417_n150# 0.43fF
C52 a_255_n150# a_159_n150# 0.43fF
C53 a_351_n150# a_255_n150# 0.43fF
C54 a_n509_n150# w_n647_n369# 0.14fF
C55 a_447_n150# VSUBS 0.03fF
C56 a_351_n150# VSUBS 0.03fF
C57 a_255_n150# VSUBS 0.03fF
C58 a_159_n150# VSUBS 0.03fF
C59 a_63_n150# VSUBS 0.03fF
C60 a_n33_n150# VSUBS 0.03fF
C61 a_n129_n150# VSUBS 0.03fF
C62 a_n225_n150# VSUBS 0.03fF
C63 a_n321_n150# VSUBS 0.03fF
C64 a_n417_n150# VSUBS 0.03fF
C65 a_n509_n150# VSUBS 0.03fF
C66 a_n465_n247# VSUBS 1.07fF
C67 w_n647_n369# VSUBS 4.87fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EDT3AT a_15_n11# a_n33_n99# w_n211_n221# a_n73_n11#
X0 a_15_n11# a_n33_n99# a_n73_n11# w_n211_n221# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_n33_n99# a_n73_n11# 0.02fF
C1 a_n33_n99# a_15_n11# 0.02fF
C2 a_15_n11# a_n73_n11# 0.15fF
C3 a_15_n11# w_n211_n221# 0.09fF
C4 a_n73_n11# w_n211_n221# 0.09fF
C5 a_n33_n99# w_n211_n221# 0.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AQR2CW a_n33_66# a_n78_n106# w_n216_n254# a_20_n106#
X0 a_20_n106# a_n33_66# a_n78_n106# w_n216_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=200000u
C0 a_20_n106# a_n78_n106# 0.21fF
C1 a_20_n106# w_n216_n254# 0.14fF
C2 a_n78_n106# w_n216_n254# 0.14fF
C3 a_n33_66# w_n216_n254# 0.12fF
.ends

.subckt sky130_fd_pr__pfet_01v8_HRYSXS VSUBS a_n33_n211# a_n78_n114# w_n216_n334#
+ a_20_n114#
X0 a_20_n114# a_n33_n211# a_n78_n114# w_n216_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=200000u
C0 a_20_n114# w_n216_n334# 0.20fF
C1 w_n216_n334# a_n78_n114# 0.20fF
C2 a_20_n114# a_n78_n114# 0.42fF
C3 a_20_n114# VSUBS 0.03fF
C4 a_n78_n114# VSUBS 0.03fF
C5 a_n33_n211# VSUBS 0.12fF
C6 w_n216_n334# VSUBS 1.66fF
.ends

.subckt inverter_csvco in vbulkn out vbulkp vdd vss
Xsky130_fd_pr__nfet_01v8_AQR2CW_0 in vss vbulkn out sky130_fd_pr__nfet_01v8_AQR2CW
Xsky130_fd_pr__pfet_01v8_HRYSXS_0 vbulkn in vdd vbulkp out sky130_fd_pr__pfet_01v8_HRYSXS
C0 in vss 0.01fF
C1 in vdd 0.01fF
C2 in out 0.11fF
C3 vdd vbulkp 0.04fF
C4 out vbulkp 0.08fF
C5 vbulkp vbulkn 2.49fF
C6 out vbulkn 0.60fF
C7 vdd vbulkn 0.06fF
C8 in vbulkn 0.54fF
C9 vss vbulkn 0.17fF
.ends

.subckt csvco_branch vctrl inverter_csvco_0/vdd in vbp cap_vco_0/t D0 out inverter_csvco_0/vss
+ vss vdd
Xsky130_fd_pr__nfet_01v8_7H8F5S_0 vctrl inverter_csvco_0/vss inverter_csvco_0/vss
+ vss vss inverter_csvco_0/vss vss vss inverter_csvco_0/vss vss inverter_csvco_0/vss
+ vss vss sky130_fd_pr__nfet_01v8_7H8F5S
Xsky130_fd_pr__pfet_01v8_8DL6ZL_0 vss inverter_csvco_0/vdd inverter_csvco_0/vdd vdd
+ inverter_csvco_0/vdd vdd vdd inverter_csvco_0/vdd vbp vdd inverter_csvco_0/vdd vdd
+ vdd vdd sky130_fd_pr__pfet_01v8_8DL6ZL
Xsky130_fd_pr__nfet_01v8_EDT3AT_0 cap_vco_0/t D0 vss out sky130_fd_pr__nfet_01v8_EDT3AT
Xinverter_csvco_0 in vss out vdd inverter_csvco_0/vdd inverter_csvco_0/vss inverter_csvco
C0 out inverter_csvco_0/vss 0.03fF
C1 D0 out 0.09fF
C2 D0 inverter_csvco_0/vss 0.02fF
C3 vdd cap_vco_0/t 0.04fF
C4 inverter_csvco_0/vss vctrl 0.87fF
C5 inverter_csvco_0/vdd cap_vco_0/t 0.10fF
C6 inverter_csvco_0/vdd in 0.01fF
C7 vdd vbp 1.21fF
C8 inverter_csvco_0/vdd vdd 1.89fF
C9 inverter_csvco_0/vdd vbp 0.75fF
C10 cap_vco_0/t out 0.70fF
C11 out in 0.06fF
C12 inverter_csvco_0/vdd out 0.02fF
C13 inverter_csvco_0/vss in 0.01fF
C14 out vss 0.93fF
C15 inverter_csvco_0/vdd vss 0.26fF
C16 in vss 0.69fF
C17 D0 vss -0.67fF
C18 vbp vss 0.13fF
C19 vdd vss 9.58fF
C20 cap_vco_0/t vss 7.22fF
C21 inverter_csvco_0/vss vss 1.79fF
C22 vctrl vss 3.06fF
.ends

.subckt ring_osc csvco_branch_0/inverter_csvco_0/vdd vctrl csvco_branch_1/inverter_csvco_0/vdd
+ csvco_branch_2/inverter_csvco_0/vdd vdd vss csvco_branch_2/vbp csvco_branch_0/inverter_csvco_0/vss
+ D0 csvco_branch_2/cap_vco_0/t out_vco
Xsky130_fd_pr__nfet_01v8_CBAU6Y_0 vss vctrl vss csvco_branch_2/vbp sky130_fd_pr__nfet_01v8_CBAU6Y
Xsky130_fd_pr__pfet_01v8_4757AC_0 vss vdd csvco_branch_2/vbp vdd csvco_branch_2/vbp
+ sky130_fd_pr__pfet_01v8_4757AC
Xcsvco_branch_0 vctrl csvco_branch_0/inverter_csvco_0/vdd out_vco csvco_branch_2/vbp
+ csvco_branch_0/cap_vco_0/t D0 csvco_branch_1/in csvco_branch_0/inverter_csvco_0/vss
+ vss vdd csvco_branch
Xcsvco_branch_2 vctrl csvco_branch_2/inverter_csvco_0/vdd csvco_branch_2/in csvco_branch_2/vbp
+ csvco_branch_2/cap_vco_0/t D0 out_vco csvco_branch_2/inverter_csvco_0/vss vss vdd
+ csvco_branch
Xcsvco_branch_1 vctrl csvco_branch_1/inverter_csvco_0/vdd csvco_branch_1/in csvco_branch_2/vbp
+ csvco_branch_1/cap_vco_0/t D0 csvco_branch_2/in csvco_branch_1/inverter_csvco_0/vss
+ vss vdd csvco_branch
C0 D0 csvco_branch_0/inverter_csvco_0/vss 0.49fF
C1 vdd csvco_branch_0/inverter_csvco_0/vdd 0.13fF
C2 csvco_branch_2/vbp csvco_branch_0/inverter_csvco_0/vss 0.06fF
C3 vdd csvco_branch_1/inverter_csvco_0/vdd 0.19fF
C4 csvco_branch_0/cap_vco_0/t out_vco 0.03fF
C5 csvco_branch_2/vbp vdd 1.49fF
C6 D0 csvco_branch_1/inverter_csvco_0/vss 0.68fF
C7 csvco_branch_2/inverter_csvco_0/vdd vdd 0.10fF
C8 vctrl D0 4.41fF
C9 csvco_branch_2/vbp csvco_branch_0/inverter_csvco_0/vdd 0.06fF
C10 D0 csvco_branch_2/inverter_csvco_0/vss 0.68fF
C11 vctrl csvco_branch_2/vbp 0.06fF
C12 csvco_branch_2/in out_vco 0.58fF
C13 csvco_branch_1/cap_vco_0/t out_vco 0.03fF
C14 csvco_branch_1/in out_vco 0.76fF
C15 csvco_branch_2/in vss 1.60fF
C16 csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C17 csvco_branch_1/cap_vco_0/t vss 7.10fF
C18 csvco_branch_1/inverter_csvco_0/vss vss 0.72fF
C19 csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C20 csvco_branch_2/cap_vco_0/t vss 7.10fF
C21 csvco_branch_2/inverter_csvco_0/vss vss 0.62fF
C22 csvco_branch_1/in vss 1.58fF
C23 csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C24 out_vco vss 0.67fF
C25 D0 vss -1.55fF
C26 vdd vss 31.40fF
C27 csvco_branch_0/cap_vco_0/t vss 7.10fF
C28 csvco_branch_0/inverter_csvco_0/vss vss 0.66fF
C29 vctrl vss 11.02fF
C30 csvco_branch_2/vbp vss 0.77fF
.ends

.subckt ring_osc_buffer vss in_vco vdd o1 out_div out_pad
Xinverter_min_x4_0 o1 vss out_div vdd inverter_min_x4
Xinverter_min_x4_1 out_div vss out_pad vdd inverter_min_x4
Xinverter_min_x2_0 in_vco o1 vss vdd inverter_min_x2
C0 vdd o1 0.09fF
C1 o1 out_div 0.11fF
C2 vdd out_div 0.17fF
C3 vdd out_pad 0.10fF
C4 out_pad out_div 0.15fF
C5 in_vco vss 0.83fF
C6 out_pad vss 0.70fF
C7 out_div vss 3.00fF
C8 vdd vss 14.54fF
C9 o1 vss 2.72fF
.ends

.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X a_194_125# a_355_368# a_455_87#
+ a_158_392#
X0 X B a_455_87# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 X a_194_125# a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_194_125# B a_158_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_158_392# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_355_368# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_194_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 a_455_87# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND B a_194_125# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X9 VGND a_194_125# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
C0 a_355_368# B 0.08fF
C1 VPWR X 0.07fF
C2 a_194_125# a_355_368# 0.51fF
C3 A B 0.28fF
C4 a_194_125# A 0.18fF
C5 VGND B 0.10fF
C6 a_194_125# VGND 0.25fF
C7 A a_355_368# 0.02fF
C8 X B 0.13fF
C9 a_194_125# X 0.29fF
C10 VGND A 0.31fF
C11 X a_355_368# 0.17fF
C12 VPWR B 0.09fF
C13 VPWR a_194_125# 0.33fF
C14 VPWR a_355_368# 0.37fF
C15 VGND X 0.28fF
C16 a_194_125# a_158_392# 0.06fF
C17 VPWR VPB 0.06fF
C18 VPWR A 0.15fF
C19 VPWR VGND 0.01fF
C20 a_194_125# B 0.57fF
C21 VGND VNB 0.78fF
C22 X VNB 0.21fF
C23 VPWR VNB 0.78fF
C24 B VNB 0.56fF
C25 A VNB 0.70fF
C26 VPB VNB 0.77fF
C27 a_355_368# VNB 0.08fF
C28 a_194_125# VNB 0.40fF
.ends

.subckt sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X a_143_136# a_56_136#
X0 VGND B a_143_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 X a_56_136# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VPWR B a_56_136# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_143_136# A a_56_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_56_136# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 X a_56_136# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
C0 a_56_136# VGND 0.06fF
C1 VGND A 0.21fF
C2 a_56_136# A 0.17fF
C3 B VPWR 0.02fF
C4 VPWR VPB 0.04fF
C5 VPWR X 0.20fF
C6 B X 0.02fF
C7 B VGND 0.03fF
C8 VGND X 0.15fF
C9 a_56_136# VPWR 0.57fF
C10 a_56_136# B 0.30fF
C11 a_56_136# X 0.26fF
C12 VPWR A 0.07fF
C13 B A 0.08fF
C14 VGND VNB 0.50fF
C15 X VNB 0.23fF
C16 VPWR VNB 0.50fF
C17 B VNB 0.24fF
C18 A VNB 0.36fF
C19 VPB VNB 0.48fF
C20 a_56_136# VNB 0.38fF
.ends

.subckt sky130_fd_sc_hs__or2_1 A B VGND VNB VPB VPWR X a_152_368# a_63_368#
X0 VPWR A a_152_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_152_368# B a_63_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 X a_63_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 X a_63_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_63_368# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X5 VGND A a_63_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
C0 VGND B 0.11fF
C1 B a_63_368# 0.14fF
C2 VGND X 0.16fF
C3 VPWR B 0.01fF
C4 a_63_368# X 0.33fF
C5 a_63_368# A 0.28fF
C6 VPWR X 0.18fF
C7 VPWR A 0.05fF
C8 a_152_368# a_63_368# 0.03fF
C9 VGND a_63_368# 0.27fF
C10 B A 0.10fF
C11 VPWR VPB 0.04fF
C12 VPWR a_63_368# 0.29fF
C13 X A 0.02fF
C14 VGND VNB 0.53fF
C15 X VNB 0.24fF
C16 A VNB 0.21fF
C17 B VNB 0.31fF
C18 VPWR VNB 0.46fF
C19 VPB VNB 0.48fF
C20 a_63_368# VNB 0.37fF
.ends

.subckt div_by_5 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in DFlipFlop_1/latch_diff_0/D
+ nCLK DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/D DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in
+ vdd DFlipFlop_2/latch_diff_0/nD Q0 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ CLK DFlipFlop_2/latch_diff_1/D vss DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ sky130_fd_sc_hs__and2_1_0/a_56_136# nQ0 DFlipFlop_1/latch_diff_1/nD CLK_5 DFlipFlop_3/latch_diff_0/nD
+ nQ2 DFlipFlop_0/latch_diff_0/D DFlipFlop_2/latch_diff_1/nD DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_1/latch_diff_1/D Q1 DFlipFlop_2/D DFlipFlop_3/latch_diff_0/D DFlipFlop_1/D
+ sky130_fd_sc_hs__xor2_1_0/a_355_368# DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ DFlipFlop_3/latch_diff_1/nD DFlipFlop_0/latch_diff_1/D Q1_shift DFlipFlop_0/latch_diff_0/nD
+ DFlipFlop_2/nQ DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop_2/latch_diff_0/D
+ sky130_fd_sc_hs__xor2_1_0/a_158_392# DFlipFlop_3/latch_diff_1/D sky130_fd_sc_hs__or2_1_0/a_63_368#
+ DFlipFlop_1/latch_diff_0/nD sky130_fd_sc_hs__and2_1_1/a_143_136# DFlipFlop_0/Q sky130_fd_sc_hs__and2_1_1/a_56_136#
+ sky130_fd_sc_hs__xor2_1_0/a_194_125# DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ sky130_fd_sc_hs__and2_1_0/a_143_136#
Xsky130_fd_sc_hs__xor2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_2/D sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ sky130_fd_sc_hs__xor2_1_0/a_355_368# sky130_fd_sc_hs__xor2_1_0/a_455_87# sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ sky130_fd_sc_hs__xor2_1
XDFlipFlop_0 DFlipFlop_0/latch_diff_0/m1_657_280# vss DFlipFlop_0/latch_diff_1/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ nQ2 DFlipFlop_0/Q DFlipFlop_0/latch_diff_1/nD DFlipFlop_0/D DFlipFlop_0/latch_diff_1/m1_657_280#
+ DFlipFlop_0/latch_diff_0/D vdd CLK DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ nCLK DFlipFlop_0/latch_diff_0/nD DFlipFlop
XDFlipFlop_1 DFlipFlop_1/latch_diff_0/m1_657_280# vss DFlipFlop_1/latch_diff_1/D DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in
+ nQ0 Q0 DFlipFlop_1/latch_diff_1/nD DFlipFlop_1/D DFlipFlop_1/latch_diff_1/m1_657_280#
+ DFlipFlop_1/latch_diff_0/D vdd CLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ nCLK DFlipFlop_1/latch_diff_0/nD DFlipFlop
XDFlipFlop_2 DFlipFlop_2/latch_diff_0/m1_657_280# vss DFlipFlop_2/latch_diff_1/D DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_2/nQ Q1 DFlipFlop_2/latch_diff_1/nD DFlipFlop_2/D DFlipFlop_2/latch_diff_1/m1_657_280#
+ DFlipFlop_2/latch_diff_0/D vdd CLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ nCLK DFlipFlop_2/latch_diff_0/nD DFlipFlop
XDFlipFlop_3 DFlipFlop_3/latch_diff_0/m1_657_280# vss DFlipFlop_3/latch_diff_1/D DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in
+ DFlipFlop_3/nQ Q1_shift DFlipFlop_3/latch_diff_1/nD Q1 DFlipFlop_3/latch_diff_1/m1_657_280#
+ DFlipFlop_3/latch_diff_0/D vdd nCLK DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out
+ CLK DFlipFlop_3/latch_diff_0/nD DFlipFlop
Xsky130_fd_sc_hs__and2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_0/D sky130_fd_sc_hs__and2_1_0/a_143_136#
+ sky130_fd_sc_hs__and2_1_0/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__and2_1_1 nQ2 nQ0 vss vss vdd vdd DFlipFlop_1/D sky130_fd_sc_hs__and2_1_1/a_143_136#
+ sky130_fd_sc_hs__and2_1_1/a_56_136# sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__or2_1_0 Q1 Q1_shift vss vss vdd vdd CLK_5 sky130_fd_sc_hs__or2_1_0/a_152_368#
+ sky130_fd_sc_hs__or2_1_0/a_63_368# sky130_fd_sc_hs__or2_1
C0 DFlipFlop_3/latch_diff_0/nD nCLK 0.08fF
C1 DFlipFlop_1/latch_diff_1/m1_657_280# nQ0 0.21fF
C2 CLK DFlipFlop_1/latch_diff_1/D 0.14fF
C3 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vdd 0.03fF
C4 DFlipFlop_1/latch_diff_1/D Q1 -0.10fF
C5 DFlipFlop_1/D sky130_fd_sc_hs__and2_1_1/a_56_136# 0.04fF
C6 DFlipFlop_1/latch_diff_1/m1_657_280# DFlipFlop_2/D 0.04fF
C7 DFlipFlop_1/latch_diff_1/m1_657_280# nCLK 0.28fF
C8 vdd sky130_fd_sc_hs__and2_1_1/a_56_136# 0.04fF
C9 DFlipFlop_2/latch_diff_1/nD nCLK 0.16fF
C10 vdd DFlipFlop_1/D 0.25fF
C11 vdd sky130_fd_sc_hs__and2_1_0/a_56_136# 0.02fF
C12 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out Q1 0.15fF
C13 DFlipFlop_1/latch_diff_1/m1_657_280# Q0 0.01fF
C14 DFlipFlop_2/nQ vdd 0.02fF
C15 CLK_5 vdd 0.15fF
C16 nCLK DFlipFlop_2/latch_diff_1/D 0.08fF
C17 CLK DFlipFlop_1/latch_diff_0/nD 0.08fF
C18 CLK sky130_fd_sc_hs__and2_1_1/a_56_136# 0.06fF
C19 CLK DFlipFlop_3/latch_diff_1/D 0.08fF
C20 DFlipFlop_0/latch_diff_1/D Q0 0.23fF
C21 CLK DFlipFlop_1/D 0.21fF
C22 CLK sky130_fd_sc_hs__and2_1_1/a_143_136# 0.03fF
C23 DFlipFlop_3/latch_diff_1/D Q1 0.79fF
C24 nCLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in -0.33fF
C25 CLK DFlipFlop_2/nQ 0.13fF
C26 Q1 DFlipFlop_1/D 0.03fF
C27 nCLK DFlipFlop_3/latch_diff_0/m1_657_280# 0.27fF
C28 Q1 sky130_fd_sc_hs__and2_1_0/a_56_136# 0.14fF
C29 Q1 DFlipFlop_2/latch_diff_0/D 0.42fF
C30 DFlipFlop_2/nQ Q1 0.31fF
C31 CLK vdd 0.41fF
C32 Q1 vdd 9.49fF
C33 CLK DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out -0.31fF
C34 vdd DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.02fF
C35 DFlipFlop_1/latch_diff_0/m1_657_280# nQ0 0.25fF
C36 DFlipFlop_2/latch_diff_1/m1_657_280# Q1 0.03fF
C37 CLK Q1 -0.10fF
C38 Q0 DFlipFlop_0/D 0.39fF
C39 sky130_fd_sc_hs__xor2_1_0/a_194_125# DFlipFlop_2/D 0.08fF
C40 nCLK sky130_fd_sc_hs__xor2_1_0/a_194_125# 0.11fF
C41 Q1 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.09fF
C42 CLK DFlipFlop_0/latch_diff_0/m1_657_280# 0.28fF
C43 sky130_fd_sc_hs__xor2_1_0/a_194_125# Q0 0.26fF
C44 Q1 DFlipFlop_0/latch_diff_0/D 0.15fF
C45 CLK DFlipFlop_0/latch_diff_1/nD 0.02fF
C46 DFlipFlop_1/latch_diff_0/D nQ0 0.09fF
C47 Q1 DFlipFlop_0/latch_diff_1/nD 0.10fF
C48 vdd DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in 0.03fF
C49 DFlipFlop_1/latch_diff_1/D nQ0 0.91fF
C50 nCLK DFlipFlop_3/nQ 0.02fF
C51 nCLK DFlipFlop_1/latch_diff_0/D 0.11fF
C52 CLK DFlipFlop_2/latch_diff_0/m1_657_280# 0.28fF
C53 CLK DFlipFlop_1/latch_diff_1/nD 0.09fF
C54 CLK DFlipFlop_3/latch_diff_1/nD 0.16fF
C55 Q1 DFlipFlop_1/latch_diff_1/nD 0.10fF
C56 Q1 DFlipFlop_3/latch_diff_1/nD 1.24fF
C57 CLK DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in 0.03fF
C58 Q0 DFlipFlop_1/latch_diff_0/D 0.42fF
C59 nCLK DFlipFlop_1/latch_diff_1/D 0.08fF
C60 DFlipFlop_1/latch_diff_1/D Q0 0.06fF
C61 Q1 sky130_fd_sc_hs__and2_1_0/a_143_136# 0.02fF
C62 Q1 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in 0.21fF
C63 DFlipFlop_1/latch_diff_0/nD nQ0 0.08fF
C64 nCLK DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out 0.05fF
C65 sky130_fd_sc_hs__and2_1_1/a_56_136# nQ0 0.01fF
C66 DFlipFlop_1/D nQ0 0.12fF
C67 sky130_fd_sc_hs__and2_1_1/a_143_136# nQ0 0.04fF
C68 Q1_shift sky130_fd_sc_hs__or2_1_0/a_63_368# -0.27fF
C69 vdd nQ0 0.11fF
C70 nCLK DFlipFlop_3/latch_diff_1/D 0.14fF
C71 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out DFlipFlop_1/D 0.03fF
C72 nCLK DFlipFlop_1/D 0.14fF
C73 nCLK DFlipFlop_2/latch_diff_0/D 0.11fF
C74 nCLK DFlipFlop_2/nQ 0.09fF
C75 nQ2 sky130_fd_sc_hs__and2_1_1/a_56_136# 0.01fF
C76 DFlipFlop_2/D vdd 0.07fF
C77 Q0 sky130_fd_sc_hs__and2_1_0/a_56_136# 0.17fF
C78 Q0 DFlipFlop_1/D 0.07fF
C79 nQ2 sky130_fd_sc_hs__and2_1_1/a_143_136# 0.01fF
C80 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vdd 0.02fF
C81 CLK nQ0 0.19fF
C82 nCLK vdd 0.34fF
C83 Q1 nQ0 0.06fF
C84 nCLK DFlipFlop_0/latch_diff_1/m1_657_280# 0.28fF
C85 nQ2 vdd 0.04fF
C86 Q0 vdd 5.33fF
C87 nCLK DFlipFlop_2/latch_diff_1/m1_657_280# 0.28fF
C88 nQ2 DFlipFlop_0/latch_diff_1/m1_657_280# 0.05fF
C89 CLK DFlipFlop_2/D 0.14fF
C90 sky130_fd_sc_hs__xor2_1_0/a_355_368# vdd 0.03fF
C91 CLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out 0.15fF
C92 Q1 DFlipFlop_2/D 0.10fF
C93 nCLK Q1 -0.01fF
C94 CLK DFlipFlop_0/Q 0.08fF
C95 Q1 DFlipFlop_0/Q 0.13fF
C96 CLK nQ2 0.17fF
C97 CLK Q0 0.08fF
C98 nQ2 Q1 0.07fF
C99 Q0 Q1 9.65fF
C100 Q0 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.33fF
C101 DFlipFlop_3/nQ Q1_shift 0.04fF
C102 nCLK DFlipFlop_0/latch_diff_1/nD 0.05fF
C103 DFlipFlop_1/latch_diff_1/nD nQ0 0.88fF
C104 Q0 DFlipFlop_0/latch_diff_0/D 0.42fF
C105 Q0 DFlipFlop_0/latch_diff_1/nD 0.21fF
C106 DFlipFlop_3/latch_diff_0/nD Q1 0.08fF
C107 nCLK DFlipFlop_1/latch_diff_1/nD 0.16fF
C108 nCLK DFlipFlop_3/latch_diff_1/nD 0.09fF
C109 Q0 DFlipFlop_1/latch_diff_1/nD 0.21fF
C110 sky130_fd_sc_hs__or2_1_0/a_152_368# Q1_shift -0.04fF
C111 nCLK DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in 0.14fF
C112 DFlipFlop_2/latch_diff_1/nD CLK 0.09fF
C113 Q0 sky130_fd_sc_hs__and2_1_0/a_143_136# 0.03fF
C114 CLK_5 sky130_fd_sc_hs__or2_1_0/a_63_368# 0.06fF
C115 vdd DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in 0.03fF
C116 DFlipFlop_2/latch_diff_1/nD Q1 0.21fF
C117 CLK DFlipFlop_3/latch_diff_1/m1_657_280# 0.27fF
C118 Q1 DFlipFlop_3/latch_diff_1/m1_657_280# 0.28fF
C119 vdd sky130_fd_sc_hs__or2_1_0/a_63_368# 0.02fF
C120 CLK DFlipFlop_2/latch_diff_1/D 0.14fF
C121 DFlipFlop_0/latch_diff_1/D CLK 0.03fF
C122 Q0 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in 0.42fF
C123 DFlipFlop_2/latch_diff_1/D Q1 0.23fF
C124 DFlipFlop_0/latch_diff_1/D Q1 0.06fF
C125 DFlipFlop_0/D sky130_fd_sc_hs__and2_1_0/a_56_136# 0.04fF
C126 vdd Q1_shift 0.10fF
C127 Q1 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in 0.20fF
C128 Q1 DFlipFlop_3/latch_diff_0/m1_657_280# 0.28fF
C129 DFlipFlop_0/D vdd 0.19fF
C130 Q1 sky130_fd_sc_hs__or2_1_0/a_63_368# 0.10fF
C131 CLK DFlipFlop_2/latch_diff_0/nD 0.08fF
C132 nCLK nQ0 0.09fF
C133 Q1 Q1_shift 0.36fF
C134 sky130_fd_sc_hs__xor2_1_0/a_194_125# vdd 0.03fF
C135 nQ2 nQ0 0.03fF
C136 Q0 nQ0 0.33fF
C137 Q1 DFlipFlop_0/D 0.13fF
C138 nCLK DFlipFlop_2/D 0.41fF
C139 DFlipFlop_0/D DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.02fF
C140 nCLK DFlipFlop_0/Q 0.11fF
C141 CLK DFlipFlop_1/latch_diff_0/m1_657_280# 0.28fF
C142 Q0 DFlipFlop_2/D 0.25fF
C143 nCLK nQ2 0.10fF
C144 nCLK Q0 0.20fF
C145 sky130_fd_sc_hs__xor2_1_0/a_455_87# DFlipFlop_2/D 0.08fF
C146 nQ2 DFlipFlop_0/Q 0.09fF
C147 nCLK sky130_fd_sc_hs__xor2_1_0/a_455_87# 0.02fF
C148 Q0 DFlipFlop_0/Q 0.21fF
C149 nQ2 Q0 0.23fF
C150 DFlipFlop_3/nQ vdd 0.02fF
C151 Q0 sky130_fd_sc_hs__xor2_1_0/a_355_368# 0.03fF
C152 CLK DFlipFlop_3/latch_diff_0/D 0.11fF
C153 Q1 DFlipFlop_3/latch_diff_0/D 0.09fF
C154 CLK DFlipFlop_3/nQ 0.01fF
C155 Q1 DFlipFlop_3/nQ 0.10fF
C156 Q1 DFlipFlop_1/latch_diff_0/D 0.18fF
C157 CLK_5 vss -0.18fF
C158 sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.38fF
C159 sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.41fF
C160 sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.38fF
C161 DFlipFlop_3/nQ vss 0.52fF
C162 Q1_shift vss -0.29fF
C163 DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.64fF
C164 DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C165 DFlipFlop_3/latch_diff_1/D vss -1.73fF
C166 DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C167 DFlipFlop_3/latch_diff_0/D vss 0.96fF
C168 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.94fF
C169 DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.85fF
C170 DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C171 DFlipFlop_2/nQ vss 0.50fF
C172 Q1 vss 8.55fF
C173 DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.72fF
C174 DFlipFlop_2/latch_diff_1/nD vss 0.58fF
C175 DFlipFlop_2/latch_diff_1/D vss -1.72fF
C176 DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C177 DFlipFlop_2/latch_diff_0/D vss 0.96fF
C178 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.89fF
C179 DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C180 DFlipFlop_2/D vss 5.34fF
C181 DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C182 nQ0 vss 3.42fF
C183 Q0 vss 0.53fF
C184 DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.62fF
C185 DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C186 DFlipFlop_1/latch_diff_1/D vss -1.73fF
C187 DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C188 DFlipFlop_1/latch_diff_0/D vss 0.96fF
C189 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C190 DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.78fF
C191 DFlipFlop_1/D vss 3.72fF
C192 DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C193 nQ2 vss 2.05fF
C194 DFlipFlop_0/Q vss -0.94fF
C195 DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.61fF
C196 nCLK vss 0.96fF
C197 DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C198 DFlipFlop_0/latch_diff_1/D vss -1.73fF
C199 DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C200 CLK vss 0.20fF
C201 DFlipFlop_0/latch_diff_0/D vss 0.96fF
C202 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.88fF
C203 DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C204 DFlipFlop_0/D vss 4.04fF
C205 DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C206 vdd vss 146.76fF
C207 sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C208 sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.42fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AZESM8 a_n63_n151# a_n33_n125# a_n255_n151# a_33_n151#
+ a_n225_n125# a_63_n125# a_n129_n125# a_n159_n151# w_n455_n335# a_225_n151# a_255_n125#
+ a_129_n151# a_159_n125# a_n317_n125#
X0 a_159_n125# a_129_n151# a_63_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n225_n125# a_n255_n151# a_n317_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_63_n125# a_33_n151# a_n33_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_n129_n125# a_n159_n151# a_n225_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n33_n125# a_n63_n151# a_n129_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_255_n125# a_225_n151# a_159_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 a_255_n125# a_63_n125# 0.13fF
C1 a_63_n125# a_n317_n125# 0.06fF
C2 a_n129_n125# a_159_n125# 0.08fF
C3 a_n225_n125# a_n317_n125# 0.36fF
C4 a_n255_n151# a_n159_n151# 0.02fF
C5 a_n159_n151# a_n63_n151# 0.02fF
C6 a_n33_n125# a_255_n125# 0.08fF
C7 a_n33_n125# a_n317_n125# 0.08fF
C8 a_n129_n125# a_63_n125# 0.13fF
C9 a_33_n151# a_129_n151# 0.02fF
C10 a_n129_n125# a_n225_n125# 0.36fF
C11 a_33_n151# a_n63_n151# 0.02fF
C12 a_159_n125# a_63_n125# 0.36fF
C13 a_n129_n125# a_n33_n125# 0.36fF
C14 a_n225_n125# a_159_n125# 0.06fF
C15 a_129_n151# a_225_n151# 0.02fF
C16 a_n129_n125# a_255_n125# 0.06fF
C17 a_n129_n125# a_n317_n125# 0.13fF
C18 a_n33_n125# a_159_n125# 0.13fF
C19 a_n225_n125# a_63_n125# 0.08fF
C20 a_255_n125# a_159_n125# 0.36fF
C21 a_n33_n125# a_63_n125# 0.36fF
C22 a_n225_n125# a_n33_n125# 0.13fF
C23 a_255_n125# w_n455_n335# 0.14fF
C24 a_159_n125# w_n455_n335# 0.08fF
C25 a_63_n125# w_n455_n335# 0.07fF
C26 a_n33_n125# w_n455_n335# 0.08fF
C27 a_n129_n125# w_n455_n335# 0.07fF
C28 a_n225_n125# w_n455_n335# 0.08fF
C29 a_n317_n125# w_n455_n335# 0.14fF
C30 a_225_n151# w_n455_n335# 0.05fF
C31 a_129_n151# w_n455_n335# 0.05fF
C32 a_33_n151# w_n455_n335# 0.05fF
C33 a_n63_n151# w_n455_n335# 0.05fF
C34 a_n159_n151# w_n455_n335# 0.05fF
C35 a_n255_n151# w_n455_n335# 0.05fF
.ends

.subckt sky130_fd_pr__pfet_01v8_XJXT7S VSUBS a_n33_n125# a_n255_n154# a_33_n154# a_n225_n125#
+ a_n159_n154# a_63_n125# a_n129_n125# a_225_n154# a_129_n154# a_255_n125# a_159_n125#
+ a_n317_n125# w_n455_n344# a_n63_n154#
X0 a_n129_n125# a_n159_n154# a_n225_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n33_n125# a_n63_n154# a_n129_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_255_n125# a_225_n154# a_159_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_159_n125# a_129_n154# a_63_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n225_n125# a_n255_n154# a_n317_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_63_n125# a_33_n154# a_n33_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
C0 w_n455_n344# a_255_n125# 0.11fF
C1 a_159_n125# a_n129_n125# 0.08fF
C2 w_n455_n344# a_n33_n125# 0.05fF
C3 a_n225_n125# a_n33_n125# 0.13fF
C4 w_n455_n344# a_63_n125# 0.04fF
C5 a_255_n125# a_n33_n125# 0.08fF
C6 a_n129_n125# a_n317_n125# 0.13fF
C7 a_n225_n125# a_63_n125# 0.08fF
C8 a_159_n125# w_n455_n344# 0.06fF
C9 a_255_n125# a_63_n125# 0.13fF
C10 a_n33_n125# a_63_n125# 0.36fF
C11 a_159_n125# a_n225_n125# 0.06fF
C12 a_n63_n154# a_n159_n154# 0.02fF
C13 a_159_n125# a_255_n125# 0.36fF
C14 w_n455_n344# a_n317_n125# 0.11fF
C15 a_159_n125# a_n33_n125# 0.13fF
C16 w_n455_n344# a_n129_n125# 0.04fF
C17 a_n225_n125# a_n317_n125# 0.36fF
C18 a_n225_n125# a_n129_n125# 0.36fF
C19 a_33_n154# a_129_n154# 0.02fF
C20 a_159_n125# a_63_n125# 0.36fF
C21 a_n129_n125# a_255_n125# 0.06fF
C22 a_n317_n125# a_n33_n125# 0.08fF
C23 a_n129_n125# a_n33_n125# 0.36fF
C24 a_33_n154# a_n63_n154# 0.02fF
C25 a_n317_n125# a_63_n125# 0.06fF
C26 a_n129_n125# a_63_n125# 0.13fF
C27 a_n255_n154# a_n159_n154# 0.02fF
C28 w_n455_n344# a_n225_n125# 0.06fF
C29 a_225_n154# a_129_n154# 0.02fF
C30 a_255_n125# VSUBS 0.03fF
C31 a_159_n125# VSUBS 0.03fF
C32 a_63_n125# VSUBS 0.03fF
C33 a_n33_n125# VSUBS 0.03fF
C34 a_n129_n125# VSUBS 0.03fF
C35 a_n225_n125# VSUBS 0.03fF
C36 a_n317_n125# VSUBS 0.03fF
C37 a_225_n154# VSUBS 0.05fF
C38 a_129_n154# VSUBS 0.05fF
C39 a_33_n154# VSUBS 0.05fF
C40 a_n63_n154# VSUBS 0.05fF
C41 a_n159_n154# VSUBS 0.05fF
C42 a_n255_n154# VSUBS 0.05fF
C43 w_n455_n344# VSUBS 2.96fF
.ends

.subckt inverter_cp_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_AZESM8_0 in vss in in vss out out in vss in out in vss out
+ sky130_fd_pr__nfet_01v8_AZESM8
Xsky130_fd_pr__pfet_01v8_XJXT7S_0 vss vdd in in vdd in out out in in out vdd out vdd
+ in sky130_fd_pr__pfet_01v8_XJXT7S
C0 out vdd 0.29fF
C1 in out 0.85fF
C2 in vdd 0.04fF
C3 vdd vss 5.90fF
C4 out vss 1.30fF
C5 in vss 1.82fF
.ends

.subckt pfd_cp_interface vss inverter_cp_x1_2/in vdd inverter_cp_x1_0/out Down QA
+ QB nDown Up nUp
Xinverter_cp_x2_0 nDown Down vss vdd inverter_cp_x2
Xinverter_cp_x2_1 Up nUp vss vdd inverter_cp_x2
Xtrans_gate_0 nDown inverter_cp_x1_0/out vss vdd trans_gate
Xinverter_cp_x1_0 inverter_cp_x1_0/out QB vss vdd inverter_cp_x1
Xinverter_cp_x1_2 Up inverter_cp_x1_2/in vss vdd inverter_cp_x1
Xinverter_cp_x1_1 inverter_cp_x1_2/in QA vss vdd inverter_cp_x1
C0 inverter_cp_x1_2/in Up 0.12fF
C1 inverter_cp_x1_2/in vdd 0.42fF
C2 inverter_cp_x1_0/out nDown 0.11fF
C3 Up vdd 0.60fF
C4 QB vdd 0.02fF
C5 Down vdd 0.09fF
C6 nUp Up 0.20fF
C7 nDown Down 0.23fF
C8 inverter_cp_x1_0/out Down 0.12fF
C9 nDown vdd 0.80fF
C10 inverter_cp_x1_0/out vdd 0.25fF
C11 nUp vdd 0.14fF
C12 QA vdd 0.02fF
C13 inverter_cp_x1_2/in vss 2.01fF
C14 QA vss 1.09fF
C15 inverter_cp_x1_0/out vss 2.00fF
C16 QB vss 1.09fF
C17 vdd vss 28.96fF
C18 nUp vss 1.32fF
C19 Up vss 2.53fF
C20 Down vss 1.26fF
C21 nDown vss 2.98fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4F35BC VSUBS a_n129_n90# w_n359_n309# a_n63_n116#
+ a_n159_n207# a_63_n90# a_n33_n90# a_n221_n90# a_159_n90#
X0 a_159_n90# a_n63_n116# a_63_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n129_n90# a_n159_n207# a_n221_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X2 a_63_n90# a_n159_n207# a_n33_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3 a_n33_n90# a_n63_n116# a_n129_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_159_n90# a_63_n90# 0.26fF
C1 w_n359_n309# a_n129_n90# 0.06fF
C2 a_n129_n90# a_n33_n90# 0.26fF
C3 a_159_n90# a_n221_n90# 0.04fF
C4 a_n221_n90# a_63_n90# 0.06fF
C5 w_n359_n309# a_n33_n90# 0.05fF
C6 a_159_n90# a_n129_n90# 0.06fF
C7 a_n129_n90# a_63_n90# 0.09fF
C8 a_159_n90# w_n359_n309# 0.09fF
C9 a_n221_n90# a_n129_n90# 0.26fF
C10 a_159_n90# a_n33_n90# 0.09fF
C11 w_n359_n309# a_63_n90# 0.06fF
C12 a_n33_n90# a_63_n90# 0.26fF
C13 a_n63_n116# a_n159_n207# 0.12fF
C14 w_n359_n309# a_n221_n90# 0.09fF
C15 a_n221_n90# a_n33_n90# 0.09fF
C16 a_159_n90# VSUBS 0.03fF
C17 a_63_n90# VSUBS 0.03fF
C18 a_n33_n90# VSUBS 0.03fF
C19 a_n129_n90# VSUBS 0.03fF
C20 a_n221_n90# VSUBS 0.03fF
C21 a_n159_n207# VSUBS 0.30fF
C22 a_n63_n116# VSUBS 0.37fF
C23 w_n359_n309# VSUBS 2.23fF
.ends

.subckt sky130_fd_pr__nfet_01v8_C3YG4M a_n33_n45# a_33_n71# a_n129_71# w_n263_n255#
+ a_n125_n45# a_63_n45#
X0 a_63_n45# a_33_n71# a_n33_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n129_71# a_n125_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_n125_n45# a_63_n45# 0.05fF
C1 a_n33_n45# a_n125_n45# 0.13fF
C2 a_n33_n45# a_63_n45# 0.13fF
C3 a_n129_71# a_33_n71# 0.04fF
C4 a_63_n45# w_n263_n255# 0.04fF
C5 a_n33_n45# w_n263_n255# 0.04fF
C6 a_n125_n45# w_n263_n255# 0.04fF
C7 a_33_n71# w_n263_n255# 0.11fF
C8 a_n129_71# w_n263_n255# 0.14fF
.ends

.subckt nor_pfd sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd A B
Xsky130_fd_pr__pfet_01v8_4F35BC_0 vss sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vdd B A sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out vdd vdd sky130_fd_pr__pfet_01v8_4F35BC
Xsky130_fd_pr__nfet_01v8_C3YG4M_0 out B A vss vss vss sky130_fd_pr__nfet_01v8_C3YG4M
C0 B A 0.24fF
C1 vdd A 0.09fF
C2 vdd sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.02fF
C3 sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# out 0.08fF
C4 A out 0.06fF
C5 sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vdd 0.02fF
C6 B out 0.40fF
C7 vdd out 0.11fF
C8 sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C9 out vss 0.45fF
C10 sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C11 A vss 0.83fF
C12 B vss 1.09fF
C13 vdd vss 3.79fF
.ends

.subckt dff_pfd vdd vss nor_pfd_2/A Q CLK nor_pfd_3/A nor_pfd_2/B Reset
Xnor_pfd_0 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_2/A nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd CLK Q nor_pfd
Xnor_pfd_1 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# Q nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd nor_pfd_2/A nor_pfd_3/A nor_pfd
Xnor_pfd_2 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_3/A nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd nor_pfd_2/A nor_pfd_2/B nor_pfd
Xnor_pfd_3 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# nor_pfd_2/B nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90#
+ vss vdd nor_pfd_3/A Reset nor_pfd
C0 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vdd 0.06fF
C1 nor_pfd_3/A nor_pfd_2/A 0.38fF
C2 vdd nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# 0.06fF
C3 vdd nor_pfd_2/A -0.01fF
C4 Q Reset 0.14fF
C5 nor_pfd_2/B Reset 0.43fF
C6 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vdd 0.06fF
C7 nor_pfd_3/A vdd 0.09fF
C8 vdd nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# 0.06fF
C9 Q nor_pfd_2/A 1.38fF
C10 nor_pfd_2/B nor_pfd_2/A 0.05fF
C11 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vdd 0.06fF
C12 nor_pfd_3/A Q 0.98fF
C13 nor_pfd_2/B nor_pfd_3/A 0.58fF
C14 Q vdd 0.08fF
C15 nor_pfd_2/B vdd 0.02fF
C16 CLK Q 0.04fF
C17 nor_pfd_3/A Reset 0.12fF
C18 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vdd 0.06fF
C19 nor_pfd_2/B Q 2.22fF
C20 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C21 nor_pfd_2/B vss 1.42fF
C22 nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C23 nor_pfd_3/A vss 3.16fF
C24 Reset vss 1.48fF
C25 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C26 nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C27 nor_pfd_2/A vss 2.56fF
C28 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C29 Q vss 2.77fF
C30 nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C31 vdd vss 16.42fF
C32 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C33 nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C34 CLK vss 0.95fF
.ends

.subckt sky130_fd_pr__nfet_01v8_ZCYAJJ w_n359_n255# a_n33_n45# a_n159_n173# a_n221_n45#
+ a_159_n45# a_n63_n71# a_n129_n45# a_63_n45#
X0 a_63_n45# a_n159_n173# a_n33_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n63_n71# a_n129_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X2 a_159_n45# a_n63_n71# a_63_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X3 a_n129_n45# a_n159_n173# a_n221_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_n129_n45# a_n221_n45# 0.13fF
C1 a_63_n45# a_n221_n45# 0.03fF
C2 a_n33_n45# a_n129_n45# 0.13fF
C3 a_63_n45# a_n33_n45# 0.13fF
C4 a_63_n45# a_n129_n45# 0.05fF
C5 a_n159_n173# a_n63_n71# 0.10fF
C6 a_159_n45# a_n221_n45# 0.02fF
C7 a_n33_n45# a_159_n45# 0.05fF
C8 a_n33_n45# a_n221_n45# 0.05fF
C9 a_159_n45# a_n129_n45# 0.03fF
C10 a_63_n45# a_159_n45# 0.13fF
C11 a_159_n45# w_n359_n255# 0.04fF
C12 a_63_n45# w_n359_n255# 0.05fF
C13 a_n33_n45# w_n359_n255# 0.05fF
C14 a_n129_n45# w_n359_n255# 0.05fF
C15 a_n221_n45# w_n359_n255# 0.08fF
C16 a_n159_n173# w_n359_n255# 0.31fF
C17 a_n63_n71# w_n359_n255# 0.31fF
.ends

.subckt sky130_fd_pr__pfet_01v8_7T83YG VSUBS a_n125_n90# a_63_n90# a_33_n187# a_n99_n187#
+ a_n33_n90# w_n263_n309#
X0 a_63_n90# a_33_n187# a_n33_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n33_n90# a_n99_n187# a_n125_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 a_n99_n187# a_33_n187# 0.04fF
C1 a_63_n90# a_n125_n90# 0.09fF
C2 a_n33_n90# a_63_n90# 0.26fF
C3 a_n33_n90# a_n125_n90# 0.26fF
C4 a_63_n90# VSUBS 0.03fF
C5 a_n33_n90# VSUBS 0.03fF
C6 a_n125_n90# VSUBS 0.03fF
C7 a_33_n187# VSUBS 0.12fF
C8 a_n99_n187# VSUBS 0.12fF
C9 w_n263_n309# VSUBS 1.21fF
.ends

.subckt sky130_fd_pr__nfet_01v8_ZXAV3F a_n73_n45# a_n33_67# a_15_n45# w_n211_n255#
X0 a_15_n45# a_n33_67# a_n73_n45# w_n211_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
C0 a_n73_n45# a_15_n45# 0.16fF
C1 a_15_n45# w_n211_n255# 0.08fF
C2 a_n73_n45# w_n211_n255# 0.06fF
C3 a_n33_67# w_n211_n255# 0.10fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4F7GBC VSUBS a_n51_n187# a_n73_n90# a_15_n90# w_n211_n309#
X0 a_15_n90# a_n51_n187# a_n73_n90# w_n211_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
C0 w_n211_n309# a_n73_n90# 0.04fF
C1 w_n211_n309# a_15_n90# 0.09fF
C2 a_15_n90# a_n73_n90# 0.31fF
C3 a_15_n90# VSUBS 0.03fF
C4 a_n73_n90# VSUBS 0.03fF
C5 a_n51_n187# VSUBS 0.12fF
C6 w_n211_n309# VSUBS 1.24fF
.ends

.subckt and_pfd a_656_410# vss out vdd A B
Xsky130_fd_pr__nfet_01v8_ZCYAJJ_0 vss a_656_410# A vss vss B sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45#
+ sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# sky130_fd_pr__nfet_01v8_ZCYAJJ
Xsky130_fd_pr__pfet_01v8_7T83YG_0 vss vdd vdd B A a_656_410# vdd sky130_fd_pr__pfet_01v8_7T83YG
Xsky130_fd_pr__nfet_01v8_ZXAV3F_0 vss a_656_410# out vss sky130_fd_pr__nfet_01v8_ZXAV3F
Xsky130_fd_pr__pfet_01v8_4F7GBC_0 vss a_656_410# vdd out vdd sky130_fd_pr__pfet_01v8_4F7GBC
C0 A a_656_410# 0.04fF
C1 A vdd 0.05fF
C2 B a_656_410# 0.30fF
C3 B sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# 0.02fF
C4 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# a_656_410# 0.07fF
C5 out a_656_410# 0.20fF
C6 out sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# 0.03fF
C7 A B 0.33fF
C8 vdd a_656_410# 0.20fF
C9 out vdd 0.10fF
C10 vdd vss 4.85fF
C11 out vss 0.47fF
C12 a_656_410# vss 1.00fF
C13 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.13fF
C14 sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.10fF
C15 A vss 0.85fF
C16 B vss 0.95fF
.ends

.subckt PFD vss vdd Down Up A B Reset
Xdff_pfd_0 vdd vss dff_pfd_0/nor_pfd_2/A Up A dff_pfd_0/nor_pfd_3/A dff_pfd_0/nor_pfd_2/B
+ Reset dff_pfd
Xdff_pfd_1 vdd vss dff_pfd_1/nor_pfd_2/A Down B dff_pfd_1/nor_pfd_3/A dff_pfd_1/nor_pfd_2/B
+ Reset dff_pfd
Xand_pfd_0 and_pfd_0/a_656_410# vss Reset vdd Up Down and_pfd
C0 Up vdd 1.62fF
C1 vdd dff_pfd_0/nor_pfd_2/A 0.13fF
C2 Down vdd 0.08fF
C3 vdd dff_pfd_1/nor_pfd_2/A 0.13fF
C4 vdd dff_pfd_0/nor_pfd_2/B 0.11fF
C5 dff_pfd_0/nor_pfd_3/A vdd 0.08fF
C6 dff_pfd_1/nor_pfd_2/B vdd 0.04fF
C7 vdd Reset 0.02fF
C8 dff_pfd_1/nor_pfd_3/A vdd 0.08fF
C9 Down Up 0.06fF
C10 and_pfd_0/a_656_410# vss 0.99fF
C11 and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C12 and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.05fF
C13 dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C14 dff_pfd_1/nor_pfd_2/B vss 1.51fF
C15 dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C16 dff_pfd_1/nor_pfd_3/A vss 3.14fF
C17 dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C18 dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C19 dff_pfd_1/nor_pfd_2/A vss 2.56fF
C20 dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C21 Down vss 3.74fF
C22 dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C23 dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C24 dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C25 B vss 1.07fF
C26 dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C27 dff_pfd_0/nor_pfd_2/B vss 1.40fF
C28 dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C29 dff_pfd_0/nor_pfd_3/A vss 3.14fF
C30 Reset vss 3.85fF
C31 dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C32 dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C33 dff_pfd_0/nor_pfd_2/A vss 2.56fF
C34 dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C35 Up vss 3.18fF
C36 dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C37 vdd vss 44.73fF
C38 dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C39 dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C40 A vss 1.07fF
.ends

.subckt top_pll_v1 vco_vctrl vdd pswitch ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd
+ charge_pump_0/w_2544_775# ring_osc_0/csvco_branch_2/vbp biasp in_ref Down vss w_13905_n238#
+ vco_D0 buffer_salida_0/a_3996_n100# ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd
+ QA charge_pump_0/w_1008_774# iref_cp ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd
+ out_to_div nDown out_to_pad Up nUp
Xloop_filter_0 lf_vc vco_vctrl vss loop_filter
Xcharge_pump_0 vss pswitch nswitch vco_vctrl vdd biasp nUp Down charge_pump_0/w_2544_775#
+ iref_cp nDown Up charge_pump_0/w_1008_774# charge_pump
Xdiv_by_2_0 vss vdd div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in out_by_2 n_out_by_2
+ out_buffer_div_2 out_to_div out_div_2 n_out_buffer_div_2 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out
+ n_out_div_2 div_by_2
Xbuffer_salida_0 buffer_salida_0/a_678_n100# out_to_pad out_to_buffer buffer_salida_0/a_3996_n100#
+ vss vdd buffer_salida
Xring_osc_0 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vco_vctrl ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd
+ ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vdd vss ring_osc_0/csvco_branch_2/vbp
+ ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vco_D0 ring_osc_0/csvco_branch_2/cap_vco_0/t
+ vco_out ring_osc
Xring_osc_buffer_0 vss vco_out vdd out_first_buffer out_to_div out_to_buffer ring_osc_buffer
Xdiv_by_5_0 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/DFlipFlop_1/latch_diff_0/D
+ n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/nD div_by_5_0/DFlipFlop_0/D div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in
+ vdd div_by_5_0/DFlipFlop_2/latch_diff_0/nD div_5_Q0 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# div_5_nQ0 div_by_5_0/DFlipFlop_1/latch_diff_1/nD
+ out_div_by_5 div_by_5_0/DFlipFlop_3/latch_diff_0/nD div_5_nQ2 div_by_5_0/DFlipFlop_0/latch_diff_0/D
+ div_by_5_0/DFlipFlop_2/latch_diff_1/nD div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_1/latch_diff_1/D div_5_Q1 div_by_5_0/DFlipFlop_2/D div_by_5_0/DFlipFlop_3/latch_diff_0/D
+ div_by_5_0/DFlipFlop_1/D div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_3/latch_diff_1/nD div_by_5_0/DFlipFlop_0/latch_diff_1/D div_5_Q1_shift
+ div_by_5_0/DFlipFlop_0/latch_diff_0/nD div_by_5_0/DFlipFlop_2/nQ div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_2/latch_diff_0/D div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ div_by_5_0/DFlipFlop_3/latch_diff_1/D div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368#
+ div_by_5_0/DFlipFlop_1/latch_diff_0/nD div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136#
+ div_by_5_0/DFlipFlop_0/Q div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136#
+ div_by_5
Xpfd_cp_interface_0 vss pfd_cp_interface_0/inverter_cp_x1_2/in vdd pfd_cp_interface_0/inverter_cp_x1_0/out
+ Down QA QB nDown Up nUp pfd_cp_interface
XPFD_0 vss vdd QB QA in_ref out_div_by_5 pfd_reset PFD
C0 div_5_Q1_shift out_div_by_5 0.05fF
C1 div_by_5_0/DFlipFlop_2/latch_diff_1/nD out_by_2 0.09fF
C2 Up pswitch 1.98fF
C3 nswitch vco_vctrl -0.06fF
C4 biasp Up 0.26fF
C5 div_by_5_0/DFlipFlop_1/latch_diff_0/nD out_by_2 0.10fF
C6 n_out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/nD 0.10fF
C7 vdd buffer_salida_0/a_678_n100# 0.24fF
C8 vdd ring_osc_0/csvco_branch_2/cap_vco_0/t 0.02fF
C9 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out out_to_div -0.12fF
C10 nUp vco_vctrl 0.02fF
C11 n_out_by_2 div_by_5_0/DFlipFlop_0/Q -0.23fF
C12 vdd nDown 0.22fF
C13 div_by_5_0/DFlipFlop_2/latch_diff_0/nD out_by_2 0.10fF
C14 vdd iref_cp 0.15fF
C15 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in out_to_div -0.16fF
C16 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# n_out_by_2 0.12fF
C17 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# out_by_2 0.10fF
C18 n_out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_0/D 0.12fF
C19 out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_1/nD 0.23fF
C20 div_by_5_0/DFlipFlop_0/Q out_by_2 0.09fF
C21 vco_vctrl div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# -0.11fF
C22 vdd QA -0.04fF
C23 vdd out_to_div 0.21fF
C24 Down nswitch 0.54fF
C25 n_out_by_2 div_5_nQ2 0.10fF
C26 n_out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/D 0.10fF
C27 nswitch nDown 0.76fF
C28 vdd vco_D0 0.03fF
C29 ring_osc_0/csvco_branch_2/vbp vco_vctrl 0.26fF
C30 n_out_by_2 vco_vctrl 0.52fF
C31 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# -0.05fF
C32 n_out_by_2 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in -0.51fF
C33 nUp nDown -0.09fF
C34 div_5_nQ2 out_by_2 0.16fF
C35 div_by_5_0/DFlipFlop_1/latch_diff_1/nD n_out_by_2 0.24fF
C36 div_by_5_0/DFlipFlop_2/latch_diff_1/D out_by_2 0.23fF
C37 div_5_Q1 out_div_by_5 0.01fF
C38 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vco_vctrl -0.36fF
C39 out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_0/nD 0.17fF
C40 vco_vctrl out_by_2 0.53fF
C41 vdd lf_vc 0.02fF
C42 vdd div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out 0.04fF
C43 div_by_5_0/DFlipFlop_1/latch_diff_1/nD out_by_2 0.09fF
C44 n_out_by_2 div_by_5_0/DFlipFlop_2/nQ 0.10fF
C45 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in out_by_2 -0.22fF
C46 Down biasp 1.24fF
C47 n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_0/D 0.24fF
C48 nDown pswitch 0.53fF
C49 div_by_5_0/DFlipFlop_2/nQ out_by_2 0.23fF
C50 biasp nDown 0.26fF
C51 vdd out_div_by_5 0.28fF
C52 vdd nUp 0.05fF
C53 n_out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_1/D 0.10fF
C54 n_out_by_2 div_5_Q1 1.04fF
C55 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out out_by_2 0.09fF
C56 div_by_5_0/DFlipFlop_0/latch_diff_1/D n_out_by_2 0.17fF
C57 vco_vctrl ring_osc_0/csvco_branch_0/inverter_csvco_0/vss 0.04fF
C58 n_out_by_2 div_by_5_0/DFlipFlop_2/D 0.19fF
C59 n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/nD 0.33fF
C60 div_by_5_0/DFlipFlop_1/latch_diff_1/D out_by_2 0.23fF
C61 div_5_Q1 out_by_2 0.42fF
C62 div_by_5_0/DFlipFlop_0/latch_diff_1/D out_by_2 0.33fF
C63 div_by_5_0/DFlipFlop_3/latch_diff_1/D n_out_by_2 0.24fF
C64 div_by_5_0/DFlipFlop_2/D out_by_2 0.22fF
C65 buffer_salida_0/a_678_n100# out_to_buffer 0.22fF
C66 n_out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_0/D 0.12fF
C67 div_by_5_0/DFlipFlop_0/latch_diff_1/nD out_by_2 0.17fF
C68 vdd Up 0.28fF
C69 n_out_by_2 div_by_5_0/DFlipFlop_1/D 0.22fF
C70 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out out_by_2 -0.04fF
C71 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392# 0.01fF
C72 out_first_buffer ring_osc_0/csvco_branch_2/cap_vco_0/t 0.03fF
C73 vdd ring_osc_0/csvco_branch_2/vbp 0.03fF
C74 vdd n_out_by_2 1.03fF
C75 n_out_by_2 div_by_5_0/DFlipFlop_3/latch_diff_0/nD 0.11fF
C76 div_5_nQ0 n_out_by_2 0.10fF
C77 div_by_5_0/DFlipFlop_3/latch_diff_1/D out_by_2 0.09fF
C78 n_out_by_2 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out -0.11fF
C79 n_out_by_2 div_by_5_0/DFlipFlop_0/D -1.48fF
C80 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136# out_by_2 -0.02fF
C81 vco_vctrl div_5_Q1 0.14fF
C82 vdd div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# 0.03fF
C83 n_out_by_2 div_5_Q0 -0.12fF
C84 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# 0.03fF
C85 div_by_5_0/DFlipFlop_1/D out_by_2 0.38fF
C86 vdd out_by_2 0.97fF
C87 out_to_buffer out_to_div 0.13fF
C88 div_5_nQ0 out_by_2 0.32fF
C89 n_out_by_2 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in 0.27fF
C90 out_by_2 div_by_5_0/DFlipFlop_0/D 0.35fF
C91 Down nDown 2.55fF
C92 iref_cp Down 0.09fF
C93 div_5_Q0 out_by_2 0.09fF
C94 div_by_5_0/DFlipFlop_3/latch_diff_0/D out_by_2 0.11fF
C95 nUp Up 2.72fF
C96 nUp pswitch 0.85fF
C97 nUp biasp -0.17fF
C98 vdd vco_vctrl -1.02fF
C99 vco_vctrl div_by_5_0/DFlipFlop_0/D -0.45fF
C100 vdd pfd_cp_interface_0/inverter_cp_x1_2/in 0.01fF
C101 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# out_div_by_5 0.18fF
C102 vdd out_to_buffer 0.07fF
C103 div_by_5_0/DFlipFlop_2/latch_diff_1/nD n_out_by_2 0.24fF
C104 vco_vctrl div_5_Q0 0.48fF
C105 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# 0.02fF
C106 n_out_by_2 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in -0.20fF
C107 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out out_by_2 0.28fF
C108 PFD_0/and_pfd_0/a_656_410# vss 0.96fF
C109 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C110 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.07fF
C111 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C112 PFD_0/dff_pfd_1/nor_pfd_2/B vss 1.40fF
C113 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C114 PFD_0/dff_pfd_1/nor_pfd_3/A vss 3.14fF
C115 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C116 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C117 PFD_0/dff_pfd_1/nor_pfd_2/A vss 2.55fF
C118 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C119 QB vss 4.46fF
C120 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C121 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C122 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C123 out_div_by_5 vss -0.40fF
C124 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C125 PFD_0/dff_pfd_0/nor_pfd_2/B vss 1.40fF
C126 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C127 PFD_0/dff_pfd_0/nor_pfd_3/A vss 3.14fF
C128 pfd_reset vss 2.17fF
C129 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C130 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C131 PFD_0/dff_pfd_0/nor_pfd_2/A vss 2.55fF
C132 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C133 QA vss 4.31fF
C134 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C135 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C136 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C137 in_ref vss 1.19fF
C138 pfd_cp_interface_0/inverter_cp_x1_2/in vss 1.85fF
C139 pfd_cp_interface_0/inverter_cp_x1_0/out vss 1.87fF
C140 nUp vss 5.50fF
C141 Up vss 2.37fF
C142 Down vss 7.92fF
C143 nDown vss -2.20fF
C144 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C145 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.38fF
C146 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.41fF
C147 div_by_5_0/DFlipFlop_3/nQ vss 0.48fF
C148 div_5_Q1_shift vss -0.14fF
C149 div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.57fF
C150 div_by_5_0/DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C151 div_by_5_0/DFlipFlop_3/latch_diff_1/D vss -1.73fF
C152 div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C153 div_by_5_0/DFlipFlop_3/latch_diff_0/D vss 0.96fF
C154 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C155 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C156 div_by_5_0/DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C157 div_by_5_0/DFlipFlop_2/nQ vss 0.48fF
C158 div_5_Q1 vss 4.28fF
C159 div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C160 div_by_5_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C161 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C162 div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C163 div_by_5_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C164 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C165 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C166 div_by_5_0/DFlipFlop_2/D vss 3.13fF
C167 div_by_5_0/DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C168 div_5_nQ0 vss 0.59fF
C169 div_5_Q0 vss 0.01fF
C170 div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C171 div_by_5_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C172 div_by_5_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C173 div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C174 div_by_5_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C175 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C176 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C177 div_by_5_0/DFlipFlop_1/D vss 3.64fF
C178 div_by_5_0/DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C179 div_5_nQ2 vss 1.24fF
C180 div_by_5_0/DFlipFlop_0/Q vss -0.94fF
C181 div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C182 n_out_by_2 vss -2.62fF
C183 div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C184 div_by_5_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C185 div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C186 out_by_2 vss -4.51fF
C187 div_by_5_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C188 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C189 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C190 div_by_5_0/DFlipFlop_0/D vss 3.96fF
C191 div_by_5_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C192 vdd vss 366.82fF
C193 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C194 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.40fF
C195 out_to_buffer vss 1.57fF
C196 out_to_div vss 4.46fF
C197 out_first_buffer vss 2.88fF
C198 ring_osc_0/csvco_branch_2/in vss 1.60fF
C199 ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C200 ring_osc_0/csvco_branch_1/cap_vco_0/t vss 7.10fF
C201 ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vss 0.52fF
C202 ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C203 ring_osc_0/csvco_branch_2/cap_vco_0/t vss 7.10fF
C204 ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vss 0.52fF
C205 ring_osc_0/csvco_branch_1/in vss 1.58fF
C206 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C207 vco_out vss 1.01fF
C208 vco_D0 vss -4.63fF
C209 ring_osc_0/csvco_branch_0/cap_vco_0/t vss 7.10fF
C210 ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vss 0.52fF
C211 ring_osc_0/csvco_branch_2/vbp vss 0.38fF
C212 out_to_pad vss 7.50fF
C213 buffer_salida_0/a_3996_n100# vss 48.29fF
C214 buffer_salida_0/a_678_n100# vss 13.38fF
C215 n_out_buffer_div_2 vss 1.63fF
C216 out_buffer_div_2 vss 1.60fF
C217 div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C218 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C219 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.89fF
C220 div_by_2_0/DFlipFlop_0/nCLK vss 1.03fF
C221 out_div_2 vss -1.30fF
C222 div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C223 div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C224 div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C225 div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C226 div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C227 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C228 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C229 n_out_div_2 vss 1.95fF
C230 div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C231 nswitch vss 3.73fF
C232 biasp vss 5.44fF
C233 iref_cp vss 2.81fF
C234 vco_vctrl vss -19.28fF
C235 pswitch vss 3.57fF
C236 lf_vc vss -59.89fF
C237 loop_filter_0/res_loop_filter_2/out vss 7.90fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_2Y8F6P VSUBS c2_n3251_n3000# m4_n3351_n3100#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
C0 m4_n3351_n3100# c2_n3251_n3000# 72.82fF
C1 m4_n3351_n3100# VSUBS 14.58fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_8P223X VSUBS a_n2017_n1317# a_n1731_n1219# a_n1879_n1219#
+ a_n2017_n61# w_n2018_n202#
X0 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X1 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X2 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X3 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X4 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X5 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X6 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X7 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X8 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X9 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X10 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X11 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X12 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X13 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X14 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X15 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X16 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X17 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X18 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X19 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X20 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X21 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X22 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X23 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X24 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X25 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X26 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X27 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X28 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X29 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X30 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X31 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X32 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X33 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X34 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X35 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X36 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X37 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X38 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X39 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X40 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X41 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X42 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X43 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X44 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X45 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X46 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X47 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X48 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X49 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
C0 w_n2018_n202# a_n2017_n61# 1.37fF
C1 w_n2018_n202# a_n1731_n1219# 19.90fF
C2 w_n2018_n202# a_n2017_n1317# 0.16fF
C3 w_n2018_n202# a_n1879_n1219# 0.25fF
C4 a_n1731_n1219# a_n2017_n61# 5.23fF
C5 a_n2017_n1317# a_n2017_n61# 2.88fF
C6 a_n1731_n1219# a_n2017_n1317# 4.73fF
C7 a_n1879_n1219# a_n2017_n61# 0.16fF
C8 a_n1879_n1219# a_n1731_n1219# 19.29fF
C9 a_n1879_n1219# a_n2017_n1317# 2.66fF
C10 a_n1879_n1219# VSUBS 1.53fF
C11 a_n2017_n1317# VSUBS 5.03fF
C12 a_n1731_n1219# VSUBS 2.60fF
C13 a_n2017_n61# VSUBS 5.10fF
C14 w_n2018_n202# VSUBS 37.43fF
.ends

.subckt bias VSUBS vdd iref_0 iref_1 iref_2 iref
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_5 VSUBS iref m1_20168_984# iref m1_20168_984#
+ vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_6 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_6/a_n1731_n1219#
+ iref_5 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_7 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219#
+ iref_6 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_9 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219#
+ iref_8 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_8 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219#
+ iref_7 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_10 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219#
+ iref_9 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_0 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_0/a_n1731_n1219#
+ iref_0 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_1 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219#
+ iref_1 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_2 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219#
+ iref_2 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_3 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219#
+ iref_3 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_4 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219#
+ iref_4 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
C0 sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219# iref_1 0.24fF
C1 iref iref_2 -0.01fF
C2 iref m1_20168_984# 0.07fF
C3 iref sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# 0.02fF
C4 vdd iref -0.07fF
C5 vdd sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219# 0.24fF
C6 iref_7 sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219# 0.24fF
C7 iref iref_1 -0.02fF
C8 iref iref_5 0.05fF
C9 iref_2 iref_3 0.05fF
C10 sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# iref_3 0.24fF
C11 vdd sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219# 0.24fF
C12 vdd sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219# 0.24fF
C13 iref iref_4 0.30fF
C14 sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# m1_20168_984# -0.39fF
C15 iref iref_8 -0.03fF
C16 sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219# iref_5 0.24fF
C17 iref_3 iref_4 0.05fF
C18 sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219# iref_8 0.24fF
C19 sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# m1_20168_984# 0.01fF
C20 vdd m1_20168_984# 0.25fF
C21 vdd sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# 0.24fF
C22 vdd sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219# 0.24fF
C23 iref_0 iref_1 0.05fF
C24 iref_2 iref_1 0.05fF
C25 iref_9 iref_8 0.05fF
C26 sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# sky130_fd_pr__pfet_01v8_lvt_8P223X_0/a_n1731_n1219# 0.67fF
C27 sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219# iref_6 0.24fF
C28 iref_7 iref_6 0.05fF
C29 iref_5 iref_6 0.05fF
C30 sky130_fd_pr__pfet_01v8_lvt_8P223X_6/a_n1731_n1219# m1_20168_984# 0.54fF
C31 iref sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# -0.15fF
C32 iref_7 iref_8 0.05fF
C33 iref_9 iref -0.01fF
C34 iref_2 sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# 0.24fF
C35 m1_20168_984# sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# 0.01fF
C36 vdd sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219# 0.24fF
C37 vdd sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# 0.24fF
C38 iref_4 VSUBS 1.17fF
C39 sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# VSUBS 2.60fF
C40 iref_3 VSUBS 0.64fF
C41 sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# VSUBS 2.60fF
C42 iref_2 VSUBS -1.26fF
C43 sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219# VSUBS 2.60fF
C44 iref_1 VSUBS -0.80fF
C45 sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# VSUBS 2.60fF
C46 iref_0 VSUBS 1.88fF
C47 iref VSUBS 32.42fF
C48 sky130_fd_pr__pfet_01v8_lvt_8P223X_0/a_n1731_n1219# VSUBS 2.60fF
C49 m1_20168_984# VSUBS 56.92fF
C50 vdd VSUBS 416.01fF
C51 iref_9 VSUBS -1.13fF
C52 sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219# VSUBS 2.60fF
C53 iref_7 VSUBS -1.38fF
C54 sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219# VSUBS 2.60fF
C55 iref_8 VSUBS -1.19fF
C56 sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219# VSUBS 2.60fF
C57 iref_6 VSUBS -1.00fF
C58 sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219# VSUBS 2.60fF
C59 iref_5 VSUBS 1.40fF
C60 sky130_fd_pr__pfet_01v8_lvt_8P223X_6/a_n1731_n1219# VSUBS 2.60fF
.ends

.subckt mimcap_decoup_1x5 VSUBS t b
Xdecap[0] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[1] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[2] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[3] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[4] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
C0 b VSUBS 68.24fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WHJTNJ VSUBS m3_n4309_50# m3_n4309_n4250# c1_n4209_n4150#
+ c1_110_n4150# m3_10_n4250#
X0 c1_n4209_n4150# m3_n4309_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 c1_110_n4150# m3_10_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2 c1_n4209_n4150# m3_n4309_50# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 c1_110_n4150# m3_10_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
C0 m3_10_n4250# c1_110_n4150# 81.11fF
C1 m3_n4309_n4250# c1_n4209_n4150# 38.10fF
C2 m3_10_n4250# m3_n4309_n4250# 1.75fF
C3 m3_n4309_50# m3_n4309_n4250# 2.63fF
C4 m3_n4309_50# c1_n4209_n4150# 38.10fF
C5 m3_n4309_50# m3_10_n4250# 1.75fF
C6 c1_110_n4150# c1_n4209_n4150# 1.32fF
C7 c1_110_n4150# VSUBS 0.12fF
C8 c1_n4209_n4150# VSUBS 0.12fF
C9 m3_n4309_n4250# VSUBS 8.68fF
C10 m3_10_n4250# VSUBS 17.92fF
C11 m3_n4309_50# VSUBS 8.68fF
.ends

.subckt cap3_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_WHJTNJ_0 VSUBS out out in in out sky130_fd_pr__cap_mim_m3_1_WHJTNJ
C0 out in 3.21fF
C1 in VSUBS -8.91fF
C2 out VSUBS 3.92fF
.ends

.subckt sky130_fd_pr__nfet_01v8_U2JGXT w_n226_n510# a_n118_n388# a_n88_n300# a_30_n300#
X0 a_30_n300# a_n118_n388# a_n88_n300# w_n226_n510# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
C0 a_n118_n388# a_n88_n300# 0.11fF
C1 a_n88_n300# a_30_n300# 0.61fF
C2 a_30_n300# w_n226_n510# 0.40fF
C3 a_n88_n300# w_n226_n510# 0.40fF
C4 a_n118_n388# w_n226_n510# 0.28fF
.ends

.subckt loop_filter_v2 vc_pex D0_cap in vss
Xcap1_loop_filter_0 vss vc_pex vss cap1_loop_filter
Xcap3_loop_filter_0 vss cap3_loop_filter_0/in vss cap3_loop_filter
Xcap2_loop_filter_0 vss in vss cap2_loop_filter
Xsky130_fd_pr__nfet_01v8_U2JGXT_0 vss D0_cap in cap3_loop_filter_0/in sky130_fd_pr__nfet_01v8_U2JGXT
Xres_loop_filter_0 vss res_loop_filter_2/out in res_loop_filter
Xres_loop_filter_1 vss res_loop_filter_2/out vc_pex res_loop_filter
Xres_loop_filter_2 vss res_loop_filter_2/out vc_pex res_loop_filter
C0 vc_pex in 0.18fF
C1 D0_cap in 0.07fF
C2 cap3_loop_filter_0/in in 0.79fF
C3 vc_pex vss -38.13fF
C4 res_loop_filter_2/out vss 8.49fF
C5 D0_cap vss 0.04fF
C6 in vss -18.54fF
C7 cap3_loop_filter_0/in vss -3.74fF
.ends

.subckt top_pll_v2 ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd pswitch vdd charge_pump_0/w_2544_775#
+ ring_osc_0/csvco_branch_2/vbp ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd in_ref
+ vco_vctrl Down w_13905_n238# vss D0_vco iref_cp ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd
+ out_to_div DO_cap nDown biasp out_to_pad Up nUp
Xcharge_pump_0 vss pswitch nswitch vco_vctrl vdd biasp nUp Down charge_pump_0/w_2544_775#
+ iref_cp nDown Up charge_pump_0/w_1008_774# charge_pump
Xloop_filter_v2_0 lf_vc DO_cap vco_vctrl vss loop_filter_v2
Xdiv_by_2_0 vss vdd div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in out_by_2 n_out_by_2
+ out_buffer_div_2 out_to_div out_div_2 n_out_buffer_div_2 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out
+ n_out_div_2 div_by_2
Xbuffer_salida_0 buffer_salida_0/a_678_n100# out_to_pad out_to_buffer buffer_salida_0/a_3996_n100#
+ vss vdd buffer_salida
Xring_osc_0 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vco_vctrl ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd
+ ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vdd vss ring_osc_0/csvco_branch_2/vbp
+ ring_osc_0/csvco_branch_0/inverter_csvco_0/vss D0_vco ring_osc_0/csvco_branch_2/cap_vco_0/t
+ vco_out ring_osc
Xring_osc_buffer_0 vss vco_out vdd out_first_buffer out_to_div out_to_buffer ring_osc_buffer
Xdiv_by_5_0 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/DFlipFlop_1/latch_diff_0/D
+ n_out_by_2 div_by_5_0/DFlipFlop_0/latch_diff_1/nD div_by_5_0/DFlipFlop_0/D div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in
+ vdd div_by_5_0/DFlipFlop_2/latch_diff_0/nD div_5_Q0 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in
+ out_by_2 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# div_5_nQ0 div_by_5_0/DFlipFlop_1/latch_diff_1/nD
+ out_div_by_5 div_by_5_0/DFlipFlop_3/latch_diff_0/nD div_5_nQ2 div_by_5_0/DFlipFlop_0/latch_diff_0/D
+ div_by_5_0/DFlipFlop_2/latch_diff_1/nD div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_1/latch_diff_1/D div_5_Q1 div_by_5_0/DFlipFlop_2/D div_by_5_0/DFlipFlop_3/latch_diff_0/D
+ div_by_5_0/DFlipFlop_1/D div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_3/latch_diff_1/nD div_by_5_0/DFlipFlop_0/latch_diff_1/D div_5_Q1_shift
+ div_by_5_0/DFlipFlop_0/latch_diff_0/nD div_by_5_0/DFlipFlop_2/nQ div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out
+ div_by_5_0/DFlipFlop_2/latch_diff_0/D div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392#
+ div_by_5_0/DFlipFlop_3/latch_diff_1/D div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368#
+ div_by_5_0/DFlipFlop_1/latch_diff_0/nD div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136#
+ div_by_5_0/DFlipFlop_0/Q div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125#
+ div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136#
+ div_by_5
Xpfd_cp_interface_0 vss pfd_cp_interface_0/inverter_cp_x1_2/in vdd pfd_cp_interface_0/inverter_cp_x1_0/out
+ Down QA QB nDown Up nUp pfd_cp_interface
XPFD_0 vss vdd QB QA in_ref out_div_by_5 pfd_reset PFD
C0 n_out_by_2 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out -0.11fF
C1 out_to_buffer out_to_div 0.13fF
C2 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# 0.03fF
C3 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_143_136# out_by_2 -0.02fF
C4 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vco_vctrl -0.36fF
C5 nswitch vco_vctrl -0.06fF
C6 div_by_5_0/DFlipFlop_3/latch_diff_0/nD n_out_by_2 0.11fF
C7 Down iref_cp 0.09fF
C8 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# vco_vctrl -0.11fF
C9 D0_vco vdd 0.03fF
C10 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# 0.12fF
C11 div_5_Q1 vco_vctrl 0.14fF
C12 nDown biasp 0.26fF
C13 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_143_136# n_out_by_2 0.02fF
C14 Down nswitch 0.54fF
C15 div_by_5_0/DFlipFlop_0/latch_diff_1/D out_by_2 0.33fF
C16 div_by_5_0/DFlipFlop_0/latch_diff_1/D n_out_by_2 0.17fF
C17 ring_osc_0/csvco_branch_2/vbp vdd 0.03fF
C18 div_5_Q1 out_by_2 0.42fF
C19 n_out_by_2 div_5_Q1 1.04fF
C20 Up biasp 0.26fF
C21 div_by_5_0/DFlipFlop_0/D vco_vctrl -0.45fF
C22 out_div_by_5 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# 0.18fF
C23 n_out_by_2 div_by_5_0/DFlipFlop_1/latch_diff_0/D 0.12fF
C24 vco_vctrl vdd -1.02fF
C25 pfd_cp_interface_0/inverter_cp_x1_2/in vdd 0.01fF
C26 div_by_5_0/DFlipFlop_0/D out_by_2 0.35fF
C27 n_out_by_2 div_by_5_0/DFlipFlop_0/D -1.48fF
C28 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in out_by_2 -0.22fF
C29 div_by_5_0/DFlipFlop_2/latch_diff_0/nD out_by_2 0.10fF
C30 ring_osc_0/csvco_branch_2/vbp vco_vctrl 0.26fF
C31 vco_vctrl ring_osc_0/csvco_branch_0/inverter_csvco_0/vss 0.04fF
C32 out_by_2 div_by_5_0/DFlipFlop_2/nQ 0.23fF
C33 n_out_by_2 div_by_5_0/DFlipFlop_2/nQ 0.10fF
C34 out_by_2 vdd 0.97fF
C35 vdd lf_vc 0.02fF
C36 div_by_5_0/DFlipFlop_0/latch_diff_1/nD out_by_2 0.17fF
C37 n_out_by_2 vdd 1.03fF
C38 div_by_5_0/DFlipFlop_1/latch_diff_1/D out_by_2 0.23fF
C39 div_by_5_0/DFlipFlop_0/latch_diff_1/nD n_out_by_2 0.33fF
C40 div_by_5_0/DFlipFlop_1/latch_diff_1/D n_out_by_2 0.10fF
C41 nUp vdd 0.05fF
C42 out_to_buffer vdd 0.07fF
C43 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out out_by_2 0.28fF
C44 nDown nswitch 0.76fF
C45 div_by_5_0/DFlipFlop_3/latch_diff_0/D out_by_2 0.11fF
C46 nUp pswitch 0.85fF
C47 vco_vctrl out_by_2 0.53fF
C48 div_5_nQ2 out_by_2 0.16fF
C49 n_out_by_2 vco_vctrl 0.52fF
C50 div_5_nQ2 n_out_by_2 0.10fF
C51 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out out_to_div -0.12fF
C52 div_by_5_0/DFlipFlop_1/latch_diff_1/nD out_by_2 0.09fF
C53 out_div_by_5 div_5_Q1 0.01fF
C54 div_by_5_0/DFlipFlop_1/latch_diff_1/nD n_out_by_2 0.24fF
C55 out_to_div div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in -0.16fF
C56 nUp vco_vctrl 0.02fF
C57 div_by_5_0/DFlipFlop_0/latch_diff_0/nD out_by_2 0.17fF
C58 out_div_by_5 div_5_Q1_shift 0.05fF
C59 div_by_5_0/DFlipFlop_3/latch_diff_1/D out_by_2 0.09fF
C60 vco_vctrl div_5_Q0 0.48fF
C61 div_by_5_0/DFlipFlop_3/latch_diff_1/D n_out_by_2 0.24fF
C62 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# out_by_2 0.10fF
C63 div_by_5_0/DFlipFlop_2/latch_diff_0/D n_out_by_2 0.12fF
C64 ring_osc_0/csvco_branch_2/cap_vco_0/t vdd 0.02fF
C65 div_5_Q0 out_by_2 0.09fF
C66 n_out_by_2 div_5_Q0 -0.12fF
C67 out_div_by_5 vdd 0.28fF
C68 nDown vdd 0.22fF
C69 div_by_5_0/DFlipFlop_0/latch_diff_0/D n_out_by_2 0.24fF
C70 Up vdd 0.28fF
C71 div_by_5_0/DFlipFlop_3/latch_diff_1/nD out_by_2 0.23fF
C72 div_by_5_0/DFlipFlop_3/latch_diff_1/nD n_out_by_2 0.10fF
C73 nDown pswitch 0.53fF
C74 out_by_2 div_by_5_0/DFlipFlop_2/D 0.22fF
C75 n_out_by_2 div_by_5_0/DFlipFlop_2/D 0.19fF
C76 div_by_5_0/DFlipFlop_0/Q out_by_2 0.09fF
C77 div_by_5_0/DFlipFlop_0/Q n_out_by_2 -0.23fF
C78 vdd buffer_salida_0/a_678_n100# 0.24fF
C79 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# n_out_by_2 -0.05fF
C80 Up pswitch 1.98fF
C81 div_by_5_0/DFlipFlop_2/latch_diff_1/nD out_by_2 0.09fF
C82 div_by_5_0/DFlipFlop_2/latch_diff_1/nD n_out_by_2 0.24fF
C83 out_by_2 div_5_nQ0 0.32fF
C84 nUp nDown -0.09fF
C85 n_out_by_2 div_5_nQ0 0.10fF
C86 n_out_by_2 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_158_392# 0.01fF
C87 nDown Down 2.55fF
C88 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in n_out_by_2 0.27fF
C89 nUp Up 2.72fF
C90 out_to_div vdd 0.21fF
C91 div_by_5_0/DFlipFlop_1/D out_by_2 0.38fF
C92 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vdd 0.04fF
C93 div_by_5_0/DFlipFlop_1/D n_out_by_2 0.22fF
C94 div_by_5_0/DFlipFlop_2/latch_diff_1/D out_by_2 0.23fF
C95 div_by_5_0/DFlipFlop_2/latch_diff_1/D n_out_by_2 0.10fF
C96 vdd iref_cp 0.15fF
C97 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in n_out_by_2 -0.20fF
C98 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in n_out_by_2 -0.51fF
C99 QA vdd -0.04fF
C100 out_to_buffer buffer_salida_0/a_678_n100# 0.22fF
C101 nUp biasp -0.17fF
C102 out_first_buffer ring_osc_0/csvco_branch_2/cap_vco_0/t 0.03fF
C103 Down biasp 1.24fF
C104 div_by_5_0/DFlipFlop_1/latch_diff_0/nD out_by_2 0.10fF
C105 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vdd 0.03fF
C106 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out out_by_2 0.09fF
C107 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out out_by_2 -0.04fF
C108 PFD_0/and_pfd_0/a_656_410# vss 0.96fF
C109 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vss 0.05fF
C110 PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vss 0.07fF
C111 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C112 PFD_0/dff_pfd_1/nor_pfd_2/B vss 1.40fF
C113 PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C114 PFD_0/dff_pfd_1/nor_pfd_3/A vss 3.14fF
C115 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C116 PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C117 PFD_0/dff_pfd_1/nor_pfd_2/A vss 2.55fF
C118 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C119 QB vss 4.46fF
C120 PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C121 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C122 PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C123 out_div_by_5 vss -0.40fF
C124 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C125 PFD_0/dff_pfd_0/nor_pfd_2/B vss 1.40fF
C126 PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C127 PFD_0/dff_pfd_0/nor_pfd_3/A vss 3.14fF
C128 pfd_reset vss 2.17fF
C129 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C130 PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C131 PFD_0/dff_pfd_0/nor_pfd_2/A vss 2.55fF
C132 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C133 QA vss 4.31fF
C134 PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C135 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vss 0.03fF
C136 PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vss 0.03fF
C137 in_ref vss 1.19fF
C138 pfd_cp_interface_0/inverter_cp_x1_2/in vss 1.85fF
C139 pfd_cp_interface_0/inverter_cp_x1_0/out vss 1.87fF
C140 nUp vss 5.50fF
C141 Up vss 2.37fF
C142 Down vss 7.92fF
C143 nDown vss -2.20fF
C144 div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vss 0.37fF
C145 div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vss 0.38fF
C146 div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vss 0.41fF
C147 div_by_5_0/DFlipFlop_3/nQ vss 0.48fF
C148 div_5_Q1_shift vss -0.14fF
C149 div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vss 0.57fF
C150 div_by_5_0/DFlipFlop_3/latch_diff_1/nD vss 0.57fF
C151 div_by_5_0/DFlipFlop_3/latch_diff_1/D vss -1.73fF
C152 div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vss 0.57fF
C153 div_by_5_0/DFlipFlop_3/latch_diff_0/D vss 0.96fF
C154 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C155 div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C156 div_by_5_0/DFlipFlop_3/latch_diff_0/nD vss 1.14fF
C157 div_by_5_0/DFlipFlop_2/nQ vss 0.48fF
C158 div_5_Q1 vss 4.28fF
C159 div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vss 0.57fF
C160 div_by_5_0/DFlipFlop_2/latch_diff_1/nD vss 0.57fF
C161 div_by_5_0/DFlipFlop_2/latch_diff_1/D vss -1.73fF
C162 div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vss 0.57fF
C163 div_by_5_0/DFlipFlop_2/latch_diff_0/D vss 0.96fF
C164 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C165 div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C166 div_by_5_0/DFlipFlop_2/D vss 3.13fF
C167 div_by_5_0/DFlipFlop_2/latch_diff_0/nD vss 1.14fF
C168 div_5_nQ0 vss 0.59fF
C169 div_5_Q0 vss 0.01fF
C170 div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vss 0.57fF
C171 div_by_5_0/DFlipFlop_1/latch_diff_1/nD vss 0.57fF
C172 div_by_5_0/DFlipFlop_1/latch_diff_1/D vss -1.73fF
C173 div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vss 0.57fF
C174 div_by_5_0/DFlipFlop_1/latch_diff_0/D vss 0.96fF
C175 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C176 div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C177 div_by_5_0/DFlipFlop_1/D vss 3.64fF
C178 div_by_5_0/DFlipFlop_1/latch_diff_0/nD vss 1.14fF
C179 div_5_nQ2 vss 1.24fF
C180 div_by_5_0/DFlipFlop_0/Q vss -0.94fF
C181 div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C182 n_out_by_2 vss -2.62fF
C183 div_by_5_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C184 div_by_5_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C185 div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C186 out_by_2 vss -4.51fF
C187 div_by_5_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C188 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C189 div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C190 div_by_5_0/DFlipFlop_0/D vss 3.96fF
C191 div_by_5_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C192 vdd vss 366.82fF
C193 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vss 0.08fF
C194 div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vss 0.40fF
C195 out_to_buffer vss 1.57fF
C196 out_to_div vss 4.46fF
C197 out_first_buffer vss 2.88fF
C198 ring_osc_0/csvco_branch_2/in vss 1.60fF
C199 ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vss 0.16fF
C200 ring_osc_0/csvco_branch_1/cap_vco_0/t vss 7.10fF
C201 ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vss 0.52fF
C202 ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vss 0.16fF
C203 ring_osc_0/csvco_branch_2/cap_vco_0/t vss 7.10fF
C204 ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vss 0.52fF
C205 ring_osc_0/csvco_branch_1/in vss 1.58fF
C206 ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vss 0.16fF
C207 vco_out vss 1.01fF
C208 D0_vco vss -4.63fF
C209 ring_osc_0/csvco_branch_0/cap_vco_0/t vss 7.10fF
C210 ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vss 0.52fF
C211 ring_osc_0/csvco_branch_2/vbp vss 0.38fF
C212 out_to_pad vss 7.50fF
C213 buffer_salida_0/a_3996_n100# vss 48.29fF
C214 buffer_salida_0/a_678_n100# vss 13.38fF
C215 n_out_buffer_div_2 vss 1.63fF
C216 out_buffer_div_2 vss 1.60fF
C217 div_by_2_0/DFlipFlop_0/CLK vss 0.31fF
C218 div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C219 div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.89fF
C220 div_by_2_0/DFlipFlop_0/nCLK vss 1.03fF
C221 out_div_2 vss -1.30fF
C222 div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vss 0.57fF
C223 div_by_2_0/DFlipFlop_0/latch_diff_1/nD vss 0.57fF
C224 div_by_2_0/DFlipFlop_0/latch_diff_1/D vss -1.73fF
C225 div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vss 0.57fF
C226 div_by_2_0/DFlipFlop_0/latch_diff_0/D vss 0.96fF
C227 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vss 1.86fF
C228 div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vss 1.76fF
C229 n_out_div_2 vss 1.95fF
C230 div_by_2_0/DFlipFlop_0/latch_diff_0/nD vss 1.14fF
C231 lf_vc vss -59.89fF
C232 loop_filter_v2_0/res_loop_filter_2/out vss 7.90fF
C233 DO_cap vss 0.01fF
C234 loop_filter_v2_0/cap3_loop_filter_0/in vss -12.03fF
C235 nswitch vss 3.73fF
C236 biasp vss 5.44fF
C237 iref_cp vss 2.81fF
C238 vco_vctrl vss -21.20fF
C239 pswitch vss 3.57fF
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[5] io_analog[7] io_analog[8] io_analog[9]
+ io_analog[4] io_analog[6] io_clamp_high[0] io_clamp_high[2] io_clamp_low[0] io_clamp_low[2]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9]
+ io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12] io_in_3v3[13] io_in_3v3[14]
+ io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18] io_in_3v3[19] io_in_3v3[1]
+ io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23] io_in_3v3[24] io_in_3v3[25]
+ io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4] io_in_3v3[5] io_in_3v3[6] io_in_3v3[7]
+ io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[2] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8]
+ io_out[9] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ user_clock2 user_irq[0] user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2
+ vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xtop_pll_v1_0 top_pll_v1_0/vco_vctrl vdda1 top_pll_v1_0/pswitch top_pll_v1_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd
+ top_pll_v1_0/charge_pump_0/w_2544_775# top_pll_v1_0/ring_osc_0/csvco_branch_2/vbp
+ top_pll_v1_0/biasp io_analog[10] top_pll_v1_0/Down vssa1 vssa1 gpio_noesd[7] top_pll_v1_0/buffer_salida_0/a_3996_n100#
+ top_pll_v1_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd top_pll_v1_0/QA top_pll_v1_0/charge_pump_0/w_1008_774#
+ bias_0/iref_2 top_pll_v1_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd top_pll_v1_0/out_to_div
+ top_pll_v1_0/nDown io_analog[9] top_pll_v1_0/Up top_pll_v1_0/nUp top_pll_v1
Xtop_pll_v1_1 top_pll_v1_1/vco_vctrl vdda1 top_pll_v1_1/pswitch top_pll_v1_1/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd
+ top_pll_v1_1/charge_pump_0/w_2544_775# top_pll_v1_1/ring_osc_0/csvco_branch_2/vbp
+ top_pll_v1_1/biasp io_analog[10] top_pll_v1_1/Down vssa1 vssa1 gpio_noesd[7] top_pll_v1_1/buffer_salida_0/a_3996_n100#
+ top_pll_v1_1/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd top_pll_v1_1/QA top_pll_v1_1/charge_pump_0/w_1008_774#
+ bias_0/iref_0 top_pll_v1_1/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd top_pll_v1_1/out_to_div
+ top_pll_v1_1/nDown io_analog[7] top_pll_v1_1/Up top_pll_v1_1/nUp top_pll_v1
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[0] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[1] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[2] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[3] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[4] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[5] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[6] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[7] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[8] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xbias_0 vssa1 vdda1 bias_0/iref_0 bias_0/iref_1 bias_0/iref_2 io_analog[5] bias
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[0] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[1] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[2] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[3] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[4] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[5] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[6] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[7] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[8] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xmimcap_decoup_1x5_0[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_0[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_0[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_1[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_1[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_1[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[0] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[1] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[2] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[3] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[4] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[5] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[6] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[7] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[8] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xmimcap_decoup_1x5_2[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_2[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_2[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_3[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_3[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_3[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_4[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_4[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_4[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_5[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_5[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_5[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xtop_pll_v2_0 top_pll_v2_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd top_pll_v2_0/pswitch
+ vdda1 top_pll_v2_0/charge_pump_0/w_2544_775# top_pll_v2_0/ring_osc_0/csvco_branch_2/vbp
+ top_pll_v2_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd io_analog[10] top_pll_v2_0/vco_vctrl
+ top_pll_v2_0/Down vssa1 vssa1 gpio_noesd[7] bias_0/iref_1 top_pll_v2_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd
+ top_pll_v2_0/out_to_div gpio_noesd[8] top_pll_v2_0/nDown top_pll_v2_0/biasp io_analog[8]
+ top_pll_v2_0/Up top_pll_v2_0/nUp top_pll_v2
C0 io_clamp_high[2] io_analog[6] 0.53fF
C1 vdda1 top_pll_v1_1/pswitch 0.48fF
C2 top_pll_v2_0/biasp vdda1 0.03fF
C3 vdda1 bias_0/iref_2 3.90fF
C4 io_analog[10] gpio_noesd[7] 29.88fF
C5 io_analog[7] top_pll_v1_1/buffer_salida_0/a_3996_n100# -0.08fF
C6 io_analog[7] bias_0/iref_2 13.22fF
C7 vdda1 gpio_noesd[7] 120.83fF
C8 top_pll_v2_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vdda1 0.17fF
C9 gpio_noesd[7] top_pll_v1_1/vco_vctrl 0.04fF
C10 vdda1 top_pll_v1_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd 0.04fF
C11 io_clamp_low[0] io_clamp_high[0] 0.53fF
C12 bias_0/iref_1 vdda1 15.26fF
C13 bias_0/iref_2 top_pll_v1_0/nDown 0.70fF
C14 io_analog[10] vdda1 0.01fF
C15 bias_0/iref_1 top_pll_v2_0/nUp 0.22fF
C16 io_analog[7] bias_0/iref_1 13.22fF
C17 io_clamp_high[0] io_analog[4] 0.53fF
C18 top_pll_v2_0/nUp vdda1 0.01fF
C19 gpio_noesd[7] top_pll_v1_0/vco_vctrl 0.05fF
C20 top_pll_v1_1/charge_pump_0/w_1008_774# bias_0/iref_0 0.21fF
C21 io_analog[7] vdda1 29.48fF
C22 vdda1 top_pll_v1_1/vco_vctrl 0.54fF
C23 top_pll_v1_0/charge_pump_0/w_2544_775# bias_0/iref_2 0.02fF
C24 bias_0/iref_1 top_pll_v2_0/nDown 0.54fF
C25 gpio_noesd[7] top_pll_v1_0/out_to_div 0.23fF
C26 vdda1 top_pll_v1_0/vco_vctrl 0.43fF
C27 top_pll_v1_1/charge_pump_0/w_2544_775# bias_0/iref_0 0.21fF
C28 vdda1 top_pll_v1_0/buffer_salida_0/a_3996_n100# 0.06fF
C29 top_pll_v1_0/ring_osc_0/csvco_branch_2/vbp vdda1 1.01fF
C30 top_pll_v1_1/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vdda1 0.12fF
C31 gpio_noesd[8] gpio_noesd[7] 1.88fF
C32 bias_0/iref_1 top_pll_v2_0/Down 0.91fF
C33 top_pll_v2_0/ring_osc_0/csvco_branch_2/vbp vdda1 2.10fF
C34 top_pll_v2_0/vco_vctrl gpio_noesd[7] 0.05fF
C35 top_pll_v1_1/Up bias_0/iref_0 0.74fF
C36 io_analog[10] gpio_noesd[8] 20.65fF
C37 vdda1 top_pll_v1_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd 0.04fF
C38 top_pll_v2_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vdda1 0.17fF
C39 io_clamp_low[2] io_analog[6] 0.53fF
C40 top_pll_v1_1/nUp bias_0/iref_0 0.74fF
C41 top_pll_v1_1/biasp bias_0/iref_0 3.13fF
C42 gpio_noesd[8] vdda1 76.96fF
C43 top_pll_v2_0/buffer_salida_0/a_3996_n100# vdda1 0.05fF
C44 top_pll_v2_0/out_to_div gpio_noesd[7] 0.23fF
C45 top_pll_v1_0/nUp bias_0/iref_2 0.70fF
C46 bias_0/iref_2 top_pll_v1_0/Down 1.11fF
C47 top_pll_v2_0/vco_vctrl vdda1 0.59fF
C48 top_pll_v2_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vdda1 0.17fF
C49 io_clamp_low[0] io_analog[4] 0.53fF
C50 top_pll_v1_1/ring_osc_0/csvco_branch_2/vbp vdda1 1.14fF
C51 bias_0/iref_1 top_pll_v2_0/charge_pump_0/w_2544_775# 0.09fF
C52 top_pll_v1_0/nUp vdda1 0.01fF
C53 vdda1 bias_0/iref_0 15.18fF
C54 top_pll_v2_0/pswitch vdda1 0.34fF
C55 vdda1 top_pll_v1_0/pswitch 0.38fF
C56 bias_0/iref_2 top_pll_v1_0/biasp 3.20fF
C57 io_analog[10] top_pll_v1_0/QA 0.03fF
C58 top_pll_v1_1/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vdda1 0.12fF
C59 io_analog[5] m3_222594_702300# 0.53fF
C60 io_analog[8] bias_0/iref_2 14.44fF
C61 io_analog[9] bias_0/iref_2 14.44fF
C62 top_pll_v1_1/out_to_div gpio_noesd[7] 0.15fF
C63 top_pll_v1_1/nDown bias_0/iref_0 0.74fF
C64 io_analog[5] m3_226242_702300# 0.53fF
C65 top_pll_v1_1/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vdda1 0.12fF
C66 top_pll_v1_1/Down bias_0/iref_0 1.08fF
C67 vdda1 top_pll_v1_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd 0.04fF
C68 vdda1 top_pll_v1_0/biasp 0.03fF
C69 bias_0/iref_1 top_pll_v2_0/Up 0.54fF
C70 io_clamp_low[2] io_clamp_high[2] 0.53fF
C71 io_analog[8] vdda1 29.93fF
C72 bias_0/iref_2 top_pll_v1_0/Up 0.70fF
C73 vdda1 io_analog[9] 30.05fF
C74 bias_0/iref_1 top_pll_v2_0/biasp 2.20fF
C75 io_in_3v3[0] vssa1 0.41fF
C76 io_oeb[26] vssa1 0.61fF
C77 io_in[0] vssa1 0.41fF
C78 io_out[26] vssa1 0.61fF
C79 io_out[0] vssa1 0.41fF
C80 io_in[26] vssa1 0.61fF
C81 io_oeb[0] vssa1 0.41fF
C82 io_in_3v3[26] vssa1 0.61fF
C83 io_in_3v3[1] vssa1 0.41fF
C84 io_oeb[25] vssa1 0.61fF
C85 io_in[1] vssa1 0.41fF
C86 io_out[25] vssa1 0.61fF
C87 io_out[1] vssa1 0.41fF
C88 io_in[25] vssa1 0.61fF
C89 io_oeb[1] vssa1 0.41fF
C90 io_in_3v3[25] vssa1 0.61fF
C91 io_in_3v3[2] vssa1 0.41fF
C92 io_oeb[24] vssa1 0.61fF
C93 io_in[2] vssa1 0.41fF
C94 io_out[24] vssa1 0.61fF
C95 io_out[2] vssa1 0.41fF
C96 io_in[24] vssa1 0.61fF
C97 io_oeb[2] vssa1 -0.20fF
C98 io_in_3v3[3] vssa1 0.41fF
C99 gpio_noesd[17] vssa1 0.61fF
C100 io_in[3] vssa1 0.41fF
C101 gpio_analog[17] vssa1 0.61fF
C102 io_out[3] vssa1 0.41fF
C103 io_oeb[3] vssa1 0.41fF
C104 io_in_3v3[4] vssa1 0.41fF
C105 io_in[4] vssa1 0.41fF
C106 io_out[4] vssa1 0.41fF
C107 io_oeb[4] vssa1 0.41fF
C108 io_oeb[23] vssa1 0.61fF
C109 io_out[23] vssa1 0.61fF
C110 io_in[23] vssa1 0.61fF
C111 io_in_3v3[23] vssa1 0.61fF
C112 gpio_noesd[16] vssa1 0.61fF
C113 io_in_3v3[5] vssa1 0.41fF
C114 io_in[5] vssa1 -0.20fF
C115 io_out[5] vssa1 0.41fF
C116 io_oeb[5] vssa1 0.41fF
C117 io_oeb[22] vssa1 0.61fF
C118 io_out[22] vssa1 0.61fF
C119 io_in[22] vssa1 0.61fF
C120 io_in_3v3[22] vssa1 0.61fF
C121 gpio_analog[15] vssa1 0.61fF
C122 io_in_3v3[6] vssa1 -0.20fF
C123 io_in[6] vssa1 0.41fF
C124 io_out[6] vssa1 0.41fF
C125 io_oeb[6] vssa1 0.41fF
C126 io_oeb[21] vssa1 0.61fF
C127 io_out[21] vssa1 0.61fF
C128 io_in[21] vssa1 0.61fF
C129 io_in_3v3[21] vssa1 0.61fF
C130 gpio_noesd[14] vssa1 0.61fF
C131 gpio_analog[14] vssa1 0.61fF
C132 vssd2 vssa1 -5.19fF
C133 vssd1 vssa1 1.13fF
C134 vdda2 vssa1 -5.19fF
C135 io_oeb[20] vssa1 0.61fF
C136 io_out[20] vssa1 0.61fF
C137 io_in[20] vssa1 0.61fF
C138 io_in_3v3[20] vssa1 0.61fF
C139 gpio_noesd[13] vssa1 0.61fF
C140 gpio_analog[13] vssa1 0.61fF
C141 gpio_analog[0] vssa1 0.41fF
C142 gpio_noesd[0] vssa1 0.41fF
C143 io_in_3v3[7] vssa1 0.41fF
C144 io_in[7] vssa1 0.41fF
C145 io_out[7] vssa1 0.41fF
C146 io_oeb[7] vssa1 0.41fF
C147 io_oeb[19] vssa1 0.61fF
C148 io_out[19] vssa1 0.61fF
C149 io_in[19] vssa1 0.61fF
C150 io_in_3v3[19] vssa1 0.61fF
C151 gpio_noesd[12] vssa1 0.61fF
C152 gpio_analog[12] vssa1 0.61fF
C153 gpio_analog[1] vssa1 0.41fF
C154 gpio_noesd[1] vssa1 0.41fF
C155 io_in_3v3[8] vssa1 0.41fF
C156 io_in[8] vssa1 0.41fF
C157 io_out[8] vssa1 -0.20fF
C158 io_oeb[8] vssa1 0.41fF
C159 io_oeb[18] vssa1 0.61fF
C160 io_out[18] vssa1 0.61fF
C161 io_in_3v3[18] vssa1 0.61fF
C162 gpio_noesd[11] vssa1 0.61fF
C163 gpio_analog[11] vssa1 0.61fF
C164 gpio_analog[2] vssa1 0.41fF
C165 gpio_noesd[2] vssa1 0.41fF
C166 io_in_3v3[9] vssa1 0.41fF
C167 io_in[9] vssa1 0.41fF
C168 io_out[9] vssa1 0.41fF
C169 io_oeb[9] vssa1 0.41fF
C170 io_oeb[17] vssa1 0.61fF
C171 io_in[17] vssa1 0.61fF
C172 io_in_3v3[17] vssa1 0.61fF
C173 gpio_noesd[10] vssa1 0.61fF
C174 gpio_analog[10] vssa1 0.61fF
C175 gpio_analog[3] vssa1 0.41fF
C176 gpio_noesd[3] vssa1 0.41fF
C177 io_in_3v3[10] vssa1 0.41fF
C178 io_in[10] vssa1 0.41fF
C179 io_out[10] vssa1 0.41fF
C180 io_oeb[10] vssa1 0.41fF
C181 io_out[16] vssa1 0.61fF
C182 io_in[16] vssa1 0.61fF
C183 io_in_3v3[16] vssa1 0.61fF
C184 gpio_noesd[9] vssa1 0.61fF
C185 gpio_analog[9] vssa1 0.61fF
C186 gpio_analog[4] vssa1 0.41fF
C187 gpio_noesd[4] vssa1 0.41fF
C188 io_in_3v3[11] vssa1 0.41fF
C189 io_in[11] vssa1 0.41fF
C190 io_out[11] vssa1 0.41fF
C191 io_oeb[11] vssa1 0.41fF
C192 io_oeb[15] vssa1 0.61fF
C193 io_out[15] vssa1 0.61fF
C194 io_in[15] vssa1 0.61fF
C195 io_in_3v3[15] vssa1 0.61fF
C196 gpio_analog[5] vssa1 0.41fF
C197 gpio_noesd[5] vssa1 0.41fF
C198 io_in_3v3[12] vssa1 0.41fF
C199 io_in[12] vssa1 0.41fF
C200 io_out[12] vssa1 0.41fF
C201 io_oeb[12] vssa1 0.41fF
C202 gpio_analog[6] vssa1 0.60fF
C203 gpio_noesd[6] vssa1 0.60fF
C204 io_in_3v3[13] vssa1 0.60fF
C205 io_in[13] vssa1 0.60fF
C206 io_out[13] vssa1 0.60fF
C207 io_oeb[13] vssa1 0.60fF
C208 vccd1 vssa1 0.85fF
C209 gpio_analog[8] vssa1 0.61fF
C210 io_oeb[14] vssa1 0.61fF
C211 io_out[14] vssa1 0.61fF
C212 io_in[14] vssa1 0.61fF
C213 io_in_3v3[14] vssa1 0.61fF
C214 io_analog[0] vssa1 -6.01fF
C215 io_analog[1] vssa1 0.76fF
C216 vssa2 vssa1 1.66fF
C217 vccd2 vssa1 0.91fF
C218 io_analog[2] vssa1 -5.85fF
C219 io_analog[3] vssa1 -5.74fF
C220 io_analog[4] vssa1 -5.03fF
C221 io_clamp_high[0] vssa1 -2.60fF
C222 io_clamp_low[0] vssa1 0.82fF
C223 io_analog[6] vssa1 -4.92fF
C224 io_clamp_high[2] vssa1 0.66fF
C225 io_clamp_low[2] vssa1 0.50fF
C226 user_irq[2] vssa1 0.63fF
C227 user_irq[1] vssa1 0.63fF
C228 user_irq[0] vssa1 0.63fF
C229 user_clock2 vssa1 0.63fF
C230 la_oenb[127] vssa1 0.63fF
C231 la_data_in[127] vssa1 0.63fF
C232 la_oenb[126] vssa1 0.63fF
C233 la_data_out[126] vssa1 0.63fF
C234 la_data_in[126] vssa1 0.63fF
C235 la_oenb[125] vssa1 0.63fF
C236 la_data_out[125] vssa1 0.63fF
C237 la_data_in[125] vssa1 0.63fF
C238 la_oenb[124] vssa1 0.63fF
C239 la_data_out[124] vssa1 0.63fF
C240 la_data_in[124] vssa1 0.63fF
C241 la_oenb[123] vssa1 0.63fF
C242 la_data_out[123] vssa1 0.63fF
C243 la_oenb[122] vssa1 0.63fF
C244 la_data_out[122] vssa1 0.63fF
C245 la_data_in[122] vssa1 0.63fF
C246 la_oenb[121] vssa1 0.63fF
C247 la_data_out[121] vssa1 0.63fF
C248 la_data_in[121] vssa1 0.63fF
C249 la_oenb[120] vssa1 0.63fF
C250 la_data_out[120] vssa1 0.63fF
C251 la_data_in[120] vssa1 0.63fF
C252 la_oenb[119] vssa1 0.63fF
C253 la_data_out[119] vssa1 0.63fF
C254 la_data_in[119] vssa1 0.63fF
C255 la_oenb[118] vssa1 0.63fF
C256 la_data_out[118] vssa1 0.63fF
C257 la_data_in[118] vssa1 0.63fF
C258 la_oenb[117] vssa1 0.63fF
C259 la_data_out[117] vssa1 0.63fF
C260 la_data_in[117] vssa1 0.63fF
C261 la_data_out[116] vssa1 0.63fF
C262 la_data_in[116] vssa1 0.63fF
C263 la_oenb[115] vssa1 0.63fF
C264 la_data_out[115] vssa1 0.63fF
C265 la_data_in[115] vssa1 0.63fF
C266 la_oenb[114] vssa1 0.63fF
C267 la_data_out[114] vssa1 0.63fF
C268 la_data_in[114] vssa1 0.63fF
C269 la_oenb[113] vssa1 0.63fF
C270 la_data_out[113] vssa1 0.63fF
C271 la_data_in[113] vssa1 0.63fF
C272 la_oenb[112] vssa1 0.63fF
C273 la_data_in[112] vssa1 0.63fF
C274 la_oenb[111] vssa1 0.63fF
C275 la_data_out[111] vssa1 0.63fF
C276 la_data_in[111] vssa1 0.63fF
C277 la_oenb[110] vssa1 0.63fF
C278 la_data_out[110] vssa1 0.63fF
C279 la_data_in[110] vssa1 0.63fF
C280 la_oenb[109] vssa1 0.63fF
C281 la_data_out[109] vssa1 0.63fF
C282 la_data_in[109] vssa1 0.63fF
C283 la_oenb[108] vssa1 0.63fF
C284 la_data_out[108] vssa1 0.63fF
C285 la_oenb[107] vssa1 0.63fF
C286 la_data_out[107] vssa1 0.63fF
C287 la_data_in[107] vssa1 0.63fF
C288 la_oenb[106] vssa1 0.63fF
C289 la_data_out[106] vssa1 0.63fF
C290 la_oenb[105] vssa1 0.63fF
C291 la_data_out[105] vssa1 0.63fF
C292 la_data_in[105] vssa1 0.63fF
C293 la_oenb[104] vssa1 0.63fF
C294 la_data_out[104] vssa1 0.63fF
C295 la_data_in[104] vssa1 0.63fF
C296 la_oenb[103] vssa1 0.63fF
C297 la_data_out[103] vssa1 0.63fF
C298 la_data_in[103] vssa1 0.63fF
C299 la_oenb[102] vssa1 0.63fF
C300 la_data_out[102] vssa1 0.63fF
C301 la_data_in[102] vssa1 0.63fF
C302 la_data_out[101] vssa1 0.63fF
C303 la_data_in[101] vssa1 0.63fF
C304 la_oenb[100] vssa1 0.63fF
C305 la_data_out[100] vssa1 0.63fF
C306 la_data_in[100] vssa1 0.63fF
C307 la_oenb[99] vssa1 0.63fF
C308 la_data_out[99] vssa1 0.63fF
C309 la_data_in[99] vssa1 0.63fF
C310 la_oenb[98] vssa1 0.63fF
C311 la_data_out[98] vssa1 0.63fF
C312 la_data_in[98] vssa1 0.63fF
C313 la_oenb[97] vssa1 0.63fF
C314 la_data_in[97] vssa1 0.63fF
C315 la_oenb[96] vssa1 0.63fF
C316 la_data_out[96] vssa1 0.63fF
C317 la_data_in[96] vssa1 0.63fF
C318 la_oenb[95] vssa1 0.63fF
C319 la_data_out[95] vssa1 0.63fF
C320 la_data_in[95] vssa1 0.63fF
C321 la_oenb[94] vssa1 0.63fF
C322 la_data_out[94] vssa1 0.63fF
C323 la_data_in[94] vssa1 0.63fF
C324 la_oenb[93] vssa1 0.63fF
C325 la_data_out[93] vssa1 0.63fF
C326 la_oenb[92] vssa1 0.63fF
C327 la_data_out[92] vssa1 0.63fF
C328 la_data_in[92] vssa1 0.63fF
C329 la_oenb[91] vssa1 0.63fF
C330 la_data_out[91] vssa1 0.63fF
C331 la_oenb[90] vssa1 0.63fF
C332 la_data_out[90] vssa1 0.63fF
C333 la_data_in[90] vssa1 0.63fF
C334 la_oenb[89] vssa1 0.63fF
C335 la_data_out[89] vssa1 0.63fF
C336 la_data_in[89] vssa1 0.63fF
C337 la_oenb[88] vssa1 0.63fF
C338 la_data_out[88] vssa1 0.63fF
C339 la_data_in[88] vssa1 0.63fF
C340 la_oenb[87] vssa1 0.63fF
C341 la_data_out[87] vssa1 0.63fF
C342 la_data_in[87] vssa1 0.63fF
C343 la_data_out[86] vssa1 0.63fF
C344 la_data_in[86] vssa1 0.63fF
C345 la_oenb[85] vssa1 0.63fF
C346 la_data_out[85] vssa1 0.63fF
C347 la_data_in[85] vssa1 0.63fF
C348 la_oenb[84] vssa1 0.63fF
C349 la_data_out[84] vssa1 0.63fF
C350 la_data_in[84] vssa1 0.63fF
C351 la_oenb[83] vssa1 0.63fF
C352 la_data_out[83] vssa1 0.63fF
C353 la_data_in[83] vssa1 0.63fF
C354 la_oenb[82] vssa1 0.63fF
C355 la_data_in[82] vssa1 0.63fF
C356 la_oenb[81] vssa1 0.63fF
C357 la_data_out[81] vssa1 0.63fF
C358 la_data_in[81] vssa1 0.63fF
C359 la_oenb[80] vssa1 0.63fF
C360 la_data_out[80] vssa1 0.63fF
C361 la_data_in[80] vssa1 0.63fF
C362 la_oenb[79] vssa1 0.63fF
C363 la_data_out[79] vssa1 0.63fF
C364 la_data_in[79] vssa1 0.63fF
C365 la_oenb[78] vssa1 0.63fF
C366 la_data_out[78] vssa1 0.63fF
C367 la_data_in[78] vssa1 0.63fF
C368 la_oenb[77] vssa1 0.63fF
C369 la_data_out[77] vssa1 0.63fF
C370 la_data_in[77] vssa1 0.63fF
C371 la_oenb[76] vssa1 0.63fF
C372 la_data_out[76] vssa1 0.63fF
C373 la_oenb[75] vssa1 0.63fF
C374 la_data_out[75] vssa1 0.63fF
C375 la_data_in[75] vssa1 0.63fF
C376 la_oenb[74] vssa1 0.63fF
C377 la_data_out[74] vssa1 0.63fF
C378 la_data_in[74] vssa1 0.63fF
C379 la_oenb[73] vssa1 0.63fF
C380 la_data_out[73] vssa1 0.63fF
C381 la_data_in[73] vssa1 0.63fF
C382 la_oenb[72] vssa1 0.63fF
C383 la_data_out[72] vssa1 0.63fF
C384 la_data_in[72] vssa1 0.63fF
C385 la_data_out[71] vssa1 0.63fF
C386 la_data_in[71] vssa1 0.63fF
C387 la_oenb[70] vssa1 0.63fF
C388 la_data_out[70] vssa1 0.63fF
C389 la_data_in[70] vssa1 0.63fF
C390 la_oenb[69] vssa1 0.63fF
C391 la_data_out[69] vssa1 0.63fF
C392 la_data_in[69] vssa1 0.63fF
C393 la_oenb[68] vssa1 0.63fF
C394 la_data_out[68] vssa1 0.63fF
C395 la_data_in[68] vssa1 0.63fF
C396 la_oenb[67] vssa1 0.63fF
C397 la_data_in[67] vssa1 0.63fF
C398 la_oenb[66] vssa1 0.63fF
C399 la_data_out[66] vssa1 0.63fF
C400 la_data_in[66] vssa1 0.63fF
C401 la_oenb[65] vssa1 0.63fF
C402 la_data_out[65] vssa1 0.26fF
C403 la_data_in[65] vssa1 0.63fF
C404 la_oenb[64] vssa1 0.63fF
C405 la_data_out[64] vssa1 0.63fF
C406 la_data_in[64] vssa1 0.63fF
C407 la_oenb[63] vssa1 0.63fF
C408 la_data_out[63] vssa1 0.63fF
C409 la_data_in[63] vssa1 0.63fF
C410 la_oenb[62] vssa1 0.63fF
C411 la_data_out[62] vssa1 0.63fF
C412 la_data_in[62] vssa1 0.63fF
C413 la_oenb[61] vssa1 0.63fF
C414 la_data_out[61] vssa1 0.63fF
C415 la_oenb[60] vssa1 0.63fF
C416 la_data_out[60] vssa1 0.63fF
C417 la_data_in[60] vssa1 0.63fF
C418 la_oenb[59] vssa1 0.63fF
C419 la_data_out[59] vssa1 0.63fF
C420 la_data_in[59] vssa1 0.63fF
C421 la_oenb[58] vssa1 0.63fF
C422 la_data_out[58] vssa1 0.63fF
C423 la_data_in[58] vssa1 0.63fF
C424 la_oenb[57] vssa1 0.63fF
C425 la_data_out[57] vssa1 0.63fF
C426 la_data_in[57] vssa1 0.63fF
C427 la_data_out[56] vssa1 0.63fF
C428 la_data_in[56] vssa1 0.63fF
C429 la_oenb[55] vssa1 0.63fF
C430 la_data_out[55] vssa1 0.63fF
C431 la_data_in[55] vssa1 0.63fF
C432 la_oenb[54] vssa1 0.63fF
C433 la_data_out[54] vssa1 0.63fF
C434 la_data_in[54] vssa1 0.63fF
C435 la_oenb[53] vssa1 0.63fF
C436 la_data_out[53] vssa1 0.63fF
C437 la_data_in[53] vssa1 0.63fF
C438 la_oenb[52] vssa1 0.63fF
C439 la_data_in[52] vssa1 0.63fF
C440 la_oenb[51] vssa1 0.63fF
C441 la_data_out[51] vssa1 0.63fF
C442 la_data_in[51] vssa1 0.63fF
C443 la_oenb[50] vssa1 0.63fF
C444 la_data_in[50] vssa1 0.63fF
C445 la_oenb[49] vssa1 0.63fF
C446 la_data_out[49] vssa1 0.63fF
C447 la_data_in[49] vssa1 0.63fF
C448 la_oenb[48] vssa1 0.63fF
C449 la_data_out[48] vssa1 0.63fF
C450 la_data_in[48] vssa1 0.63fF
C451 la_oenb[47] vssa1 0.63fF
C452 la_data_out[47] vssa1 0.63fF
C453 la_data_in[47] vssa1 0.63fF
C454 la_oenb[46] vssa1 0.63fF
C455 la_data_out[46] vssa1 0.63fF
C456 la_oenb[45] vssa1 0.63fF
C457 la_data_out[45] vssa1 0.63fF
C458 la_data_in[45] vssa1 0.63fF
C459 la_oenb[44] vssa1 0.63fF
C460 la_data_out[44] vssa1 0.63fF
C461 la_data_in[44] vssa1 0.63fF
C462 la_oenb[43] vssa1 0.63fF
C463 la_data_out[43] vssa1 0.63fF
C464 la_data_in[43] vssa1 0.63fF
C465 la_oenb[42] vssa1 0.63fF
C466 la_data_out[42] vssa1 0.63fF
C467 la_data_in[42] vssa1 0.63fF
C468 la_data_out[41] vssa1 0.63fF
C469 la_data_in[41] vssa1 0.63fF
C470 la_oenb[40] vssa1 0.63fF
C471 la_data_out[40] vssa1 0.63fF
C472 la_data_in[40] vssa1 0.63fF
C473 la_oenb[39] vssa1 0.63fF
C474 la_data_out[39] vssa1 0.63fF
C475 la_data_in[39] vssa1 0.63fF
C476 la_oenb[38] vssa1 0.63fF
C477 la_data_out[38] vssa1 0.63fF
C478 la_data_in[38] vssa1 0.63fF
C479 la_oenb[37] vssa1 0.63fF
C480 la_data_out[37] vssa1 0.26fF
C481 la_data_in[37] vssa1 0.63fF
C482 la_oenb[36] vssa1 0.63fF
C483 la_data_out[36] vssa1 0.63fF
C484 la_data_in[36] vssa1 0.63fF
C485 la_oenb[35] vssa1 0.63fF
C486 la_data_in[35] vssa1 0.63fF
C487 la_oenb[34] vssa1 0.63fF
C488 la_data_out[34] vssa1 0.63fF
C489 la_data_in[34] vssa1 0.63fF
C490 la_oenb[33] vssa1 0.63fF
C491 la_data_out[33] vssa1 0.63fF
C492 la_data_in[33] vssa1 0.63fF
C493 la_oenb[32] vssa1 0.63fF
C494 la_data_out[32] vssa1 0.63fF
C495 la_data_in[32] vssa1 0.63fF
C496 la_oenb[31] vssa1 0.63fF
C497 la_data_out[31] vssa1 0.63fF
C498 la_oenb[30] vssa1 0.63fF
C499 la_data_out[30] vssa1 0.63fF
C500 la_data_in[30] vssa1 0.63fF
C501 la_oenb[29] vssa1 0.63fF
C502 la_data_out[29] vssa1 0.63fF
C503 la_data_in[29] vssa1 0.63fF
C504 la_oenb[28] vssa1 0.63fF
C505 la_data_out[28] vssa1 0.63fF
C506 la_data_in[28] vssa1 0.63fF
C507 la_oenb[27] vssa1 0.63fF
C508 la_data_out[27] vssa1 0.63fF
C509 la_data_in[27] vssa1 0.63fF
C510 la_data_out[26] vssa1 0.63fF
C511 la_data_in[26] vssa1 0.63fF
C512 la_oenb[25] vssa1 0.63fF
C513 la_data_out[25] vssa1 0.63fF
C514 la_data_in[25] vssa1 0.63fF
C515 la_oenb[24] vssa1 0.63fF
C516 la_data_out[24] vssa1 0.63fF
C517 la_data_in[24] vssa1 0.63fF
C518 la_oenb[23] vssa1 0.63fF
C519 la_data_out[23] vssa1 0.63fF
C520 la_data_in[23] vssa1 0.63fF
C521 la_oenb[22] vssa1 0.63fF
C522 la_data_out[22] vssa1 0.63fF
C523 la_data_in[22] vssa1 0.63fF
C524 la_oenb[21] vssa1 0.63fF
C525 la_data_out[21] vssa1 0.63fF
C526 la_data_in[21] vssa1 0.63fF
C527 la_oenb[20] vssa1 0.63fF
C528 la_data_in[20] vssa1 0.63fF
C529 la_oenb[19] vssa1 0.63fF
C530 la_data_out[19] vssa1 0.63fF
C531 la_data_in[19] vssa1 0.63fF
C532 la_oenb[18] vssa1 0.63fF
C533 la_data_out[18] vssa1 0.63fF
C534 la_data_in[18] vssa1 0.63fF
C535 la_oenb[17] vssa1 0.63fF
C536 la_data_out[17] vssa1 0.63fF
C537 la_data_in[17] vssa1 0.63fF
C538 la_oenb[16] vssa1 0.63fF
C539 la_data_out[16] vssa1 0.63fF
C540 la_oenb[15] vssa1 0.63fF
C541 la_data_out[15] vssa1 0.63fF
C542 la_data_in[15] vssa1 0.63fF
C543 la_oenb[14] vssa1 0.63fF
C544 la_data_out[14] vssa1 0.63fF
C545 la_data_in[14] vssa1 0.63fF
C546 la_oenb[13] vssa1 0.63fF
C547 la_data_out[13] vssa1 0.63fF
C548 la_data_in[13] vssa1 0.63fF
C549 la_oenb[12] vssa1 0.63fF
C550 la_data_out[12] vssa1 0.63fF
C551 la_data_in[12] vssa1 0.63fF
C552 la_data_out[11] vssa1 0.63fF
C553 la_data_in[11] vssa1 0.63fF
C554 la_oenb[10] vssa1 0.63fF
C555 la_data_out[10] vssa1 0.63fF
C556 la_data_in[10] vssa1 0.63fF
C557 la_data_out[9] vssa1 0.63fF
C558 la_data_in[9] vssa1 0.63fF
C559 la_oenb[8] vssa1 0.63fF
C560 la_data_out[8] vssa1 0.63fF
C561 la_data_in[8] vssa1 0.63fF
C562 la_oenb[7] vssa1 0.63fF
C563 la_data_out[7] vssa1 0.63fF
C564 la_data_in[7] vssa1 0.63fF
C565 la_oenb[6] vssa1 0.63fF
C566 la_data_out[6] vssa1 0.63fF
C567 la_data_in[6] vssa1 0.63fF
C568 la_oenb[5] vssa1 0.63fF
C569 la_data_in[5] vssa1 0.63fF
C570 la_oenb[4] vssa1 0.63fF
C571 la_data_out[4] vssa1 0.63fF
C572 la_data_in[4] vssa1 0.63fF
C573 la_oenb[3] vssa1 0.63fF
C574 la_data_out[3] vssa1 0.63fF
C575 la_data_in[3] vssa1 0.63fF
C576 la_oenb[2] vssa1 0.63fF
C577 la_data_out[2] vssa1 0.63fF
C578 la_data_in[2] vssa1 0.63fF
C579 la_oenb[1] vssa1 0.63fF
C580 la_data_out[1] vssa1 0.63fF
C581 la_oenb[0] vssa1 0.63fF
C582 la_data_out[0] vssa1 0.63fF
C583 la_data_in[0] vssa1 0.63fF
C584 wbs_dat_o[31] vssa1 0.63fF
C585 wbs_dat_i[31] vssa1 0.63fF
C586 wbs_adr_i[31] vssa1 0.63fF
C587 wbs_dat_o[30] vssa1 0.63fF
C588 wbs_dat_i[30] vssa1 0.63fF
C589 wbs_adr_i[30] vssa1 0.63fF
C590 wbs_dat_o[29] vssa1 0.63fF
C591 wbs_dat_i[29] vssa1 0.63fF
C592 wbs_adr_i[29] vssa1 0.63fF
C593 wbs_dat_i[28] vssa1 0.63fF
C594 wbs_adr_i[28] vssa1 0.63fF
C595 wbs_dat_o[27] vssa1 0.63fF
C596 wbs_dat_i[27] vssa1 0.63fF
C597 wbs_adr_i[27] vssa1 0.63fF
C598 wbs_dat_i[26] vssa1 0.63fF
C599 wbs_adr_i[26] vssa1 0.63fF
C600 wbs_dat_o[25] vssa1 0.63fF
C601 wbs_dat_i[25] vssa1 0.63fF
C602 wbs_adr_i[25] vssa1 0.63fF
C603 wbs_dat_o[24] vssa1 0.63fF
C604 wbs_dat_i[24] vssa1 0.63fF
C605 wbs_adr_i[24] vssa1 0.63fF
C606 wbs_dat_o[23] vssa1 0.63fF
C607 wbs_dat_i[23] vssa1 0.63fF
C608 wbs_adr_i[23] vssa1 0.63fF
C609 wbs_dat_o[22] vssa1 0.63fF
C610 wbs_adr_i[22] vssa1 0.63fF
C611 wbs_dat_o[21] vssa1 0.63fF
C612 wbs_dat_i[21] vssa1 0.63fF
C613 wbs_adr_i[21] vssa1 0.63fF
C614 wbs_dat_o[20] vssa1 0.63fF
C615 wbs_dat_i[20] vssa1 0.63fF
C616 wbs_adr_i[20] vssa1 0.63fF
C617 wbs_dat_o[19] vssa1 0.63fF
C618 wbs_dat_i[19] vssa1 0.63fF
C619 wbs_adr_i[19] vssa1 0.63fF
C620 wbs_dat_o[18] vssa1 0.63fF
C621 wbs_dat_i[18] vssa1 0.63fF
C622 wbs_dat_o[17] vssa1 0.63fF
C623 wbs_dat_i[17] vssa1 0.63fF
C624 wbs_adr_i[17] vssa1 0.63fF
C625 wbs_dat_o[16] vssa1 0.63fF
C626 wbs_dat_i[16] vssa1 0.63fF
C627 wbs_adr_i[16] vssa1 0.63fF
C628 wbs_dat_o[15] vssa1 0.63fF
C629 wbs_dat_i[15] vssa1 0.63fF
C630 wbs_adr_i[15] vssa1 0.63fF
C631 wbs_dat_o[14] vssa1 0.63fF
C632 wbs_dat_i[14] vssa1 0.63fF
C633 wbs_adr_i[14] vssa1 0.63fF
C634 wbs_dat_o[13] vssa1 0.63fF
C635 wbs_dat_i[13] vssa1 0.63fF
C636 wbs_adr_i[13] vssa1 0.63fF
C637 wbs_dat_o[12] vssa1 0.63fF
C638 wbs_dat_i[12] vssa1 0.63fF
C639 wbs_adr_i[12] vssa1 0.63fF
C640 wbs_dat_i[11] vssa1 0.63fF
C641 wbs_adr_i[11] vssa1 0.63fF
C642 wbs_dat_o[10] vssa1 0.63fF
C643 wbs_dat_i[10] vssa1 0.63fF
C644 wbs_adr_i[10] vssa1 0.63fF
C645 wbs_dat_o[9] vssa1 0.63fF
C646 wbs_dat_i[9] vssa1 0.63fF
C647 wbs_adr_i[9] vssa1 0.63fF
C648 wbs_dat_o[8] vssa1 0.63fF
C649 wbs_dat_i[8] vssa1 0.63fF
C650 wbs_adr_i[8] vssa1 0.63fF
C651 wbs_dat_o[7] vssa1 0.63fF
C652 wbs_adr_i[7] vssa1 0.63fF
C653 wbs_dat_o[6] vssa1 0.63fF
C654 wbs_dat_i[6] vssa1 0.63fF
C655 wbs_adr_i[6] vssa1 0.63fF
C656 wbs_dat_o[5] vssa1 0.63fF
C657 wbs_dat_i[5] vssa1 0.63fF
C658 wbs_adr_i[5] vssa1 0.63fF
C659 wbs_dat_o[4] vssa1 0.63fF
C660 wbs_dat_i[4] vssa1 0.63fF
C661 wbs_adr_i[4] vssa1 0.63fF
C662 wbs_sel_i[3] vssa1 0.63fF
C663 wbs_dat_o[3] vssa1 0.63fF
C664 wbs_adr_i[3] vssa1 0.63fF
C665 wbs_sel_i[2] vssa1 0.63fF
C666 wbs_dat_o[2] vssa1 0.63fF
C667 wbs_dat_i[2] vssa1 0.63fF
C668 wbs_adr_i[2] vssa1 0.63fF
C669 wbs_dat_o[1] vssa1 0.63fF
C670 wbs_dat_i[1] vssa1 0.63fF
C671 wbs_adr_i[1] vssa1 0.63fF
C672 wbs_sel_i[0] vssa1 0.63fF
C673 wbs_dat_o[0] vssa1 0.63fF
C674 wbs_dat_i[0] vssa1 0.63fF
C675 wbs_adr_i[0] vssa1 0.63fF
C676 wbs_we_i vssa1 0.63fF
C677 wbs_stb_i vssa1 0.63fF
C678 wbs_cyc_i vssa1 0.63fF
C679 wbs_ack_o vssa1 0.63fF
C680 wb_rst_i vssa1 0.63fF
C681 m3_226242_702300# vssa1 -1.31fF $ **FLOATING
C682 m3_222594_702300# vssa1 0.55fF $ **FLOATING
C683 top_pll_v2_0/PFD_0/and_pfd_0/a_656_410# vssa1 0.96fF
C684 top_pll_v2_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vssa1 0.05fF
C685 top_pll_v2_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vssa1 0.05fF
C686 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C687 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_2/B vssa1 1.40fF
C688 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C689 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_3/A vssa1 3.14fF
C690 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C691 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C692 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_2/A vssa1 2.55fF
C693 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C694 top_pll_v2_0/QB vssa1 4.35fF
C695 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C696 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C697 top_pll_v2_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C698 top_pll_v2_0/out_div_by_5 vssa1 -0.40fF
C699 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C700 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_2/B vssa1 1.40fF
C701 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C702 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_3/A vssa1 3.14fF
C703 top_pll_v2_0/pfd_reset vssa1 2.17fF
C704 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C705 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C706 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_2/A vssa1 2.55fF
C707 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C708 top_pll_v2_0/QA vssa1 4.22fF
C709 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C710 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C711 top_pll_v2_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C712 top_pll_v2_0/pfd_cp_interface_0/inverter_cp_x1_2/in vssa1 1.85fF
C713 top_pll_v2_0/pfd_cp_interface_0/inverter_cp_x1_0/out vssa1 1.77fF
C714 top_pll_v2_0/nUp vssa1 5.39fF
C715 top_pll_v2_0/Up vssa1 1.85fF
C716 top_pll_v2_0/Down vssa1 6.19fF
C717 top_pll_v2_0/nDown vssa1 -3.53fF
C718 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vssa1 0.37fF
C719 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vssa1 0.38fF
C720 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vssa1 0.38fF
C721 top_pll_v2_0/div_by_5_0/DFlipFlop_3/nQ vssa1 0.48fF
C722 top_pll_v2_0/div_5_Q1_shift vssa1 -0.14fF
C723 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vssa1 0.57fF
C724 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_1/nD vssa1 0.57fF
C725 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_1/D vssa1 -1.73fF
C726 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vssa1 0.57fF
C727 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_0/D vssa1 0.96fF
C728 top_pll_v2_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C729 top_pll_v2_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C730 top_pll_v2_0/div_by_5_0/DFlipFlop_3/latch_diff_0/nD vssa1 1.14fF
C731 top_pll_v2_0/div_by_5_0/DFlipFlop_2/nQ vssa1 0.48fF
C732 top_pll_v2_0/div_5_Q1 vssa1 4.25fF
C733 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vssa1 0.57fF
C734 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD vssa1 0.57fF
C735 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D vssa1 -1.73fF
C736 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vssa1 0.57fF
C737 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D vssa1 0.96fF
C738 top_pll_v2_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C739 top_pll_v2_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C740 top_pll_v2_0/div_by_5_0/DFlipFlop_2/D vssa1 3.13fF
C741 top_pll_v2_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD vssa1 1.14fF
C742 top_pll_v2_0/div_5_nQ0 vssa1 0.59fF
C743 top_pll_v2_0/div_5_Q0 vssa1 0.01fF
C744 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vssa1 0.57fF
C745 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_1/nD vssa1 0.57fF
C746 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_1/D vssa1 -1.73fF
C747 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vssa1 0.57fF
C748 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_0/D vssa1 0.96fF
C749 top_pll_v2_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C750 top_pll_v2_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C751 top_pll_v2_0/div_by_5_0/DFlipFlop_1/D vssa1 3.64fF
C752 top_pll_v2_0/div_by_5_0/DFlipFlop_1/latch_diff_0/nD vssa1 1.14fF
C753 top_pll_v2_0/div_5_nQ2 vssa1 1.24fF
C754 top_pll_v2_0/div_by_5_0/DFlipFlop_0/Q vssa1 -0.94fF
C755 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C756 top_pll_v2_0/n_out_by_2 vssa1 -2.75fF
C757 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C758 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C759 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C760 top_pll_v2_0/out_by_2 vssa1 -5.01fF
C761 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C762 top_pll_v2_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C763 top_pll_v2_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C764 top_pll_v2_0/div_by_5_0/DFlipFlop_0/D vssa1 3.96fF
C765 top_pll_v2_0/div_by_5_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C766 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vssa1 0.08fF
C767 top_pll_v2_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vssa1 0.40fF
C768 top_pll_v2_0/out_to_buffer vssa1 1.54fF
C769 top_pll_v2_0/out_to_div vssa1 4.23fF
C770 top_pll_v2_0/out_first_buffer vssa1 2.88fF
C771 top_pll_v2_0/ring_osc_0/csvco_branch_2/in vssa1 1.60fF
C772 top_pll_v2_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vssa1 0.16fF
C773 top_pll_v2_0/ring_osc_0/csvco_branch_1/cap_vco_0/t vssa1 7.10fF
C774 top_pll_v2_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vssa1 0.52fF
C775 top_pll_v2_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vssa1 0.16fF
C776 top_pll_v2_0/ring_osc_0/csvco_branch_2/cap_vco_0/t vssa1 7.10fF
C777 top_pll_v2_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vssa1 0.52fF
C778 top_pll_v2_0/ring_osc_0/csvco_branch_1/in vssa1 1.58fF
C779 top_pll_v2_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vssa1 0.16fF
C780 top_pll_v2_0/vco_out vssa1 1.01fF
C781 top_pll_v2_0/ring_osc_0/csvco_branch_0/cap_vco_0/t vssa1 7.10fF
C782 top_pll_v2_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vssa1 0.52fF
C783 top_pll_v2_0/ring_osc_0/csvco_branch_2/vbp vssa1 0.36fF
C784 io_analog[8] vssa1 13.78fF
C785 top_pll_v2_0/buffer_salida_0/a_3996_n100# vssa1 48.23fF
C786 top_pll_v2_0/buffer_salida_0/a_678_n100# vssa1 13.21fF
C787 top_pll_v2_0/n_out_buffer_div_2 vssa1 1.63fF
C788 top_pll_v2_0/out_buffer_div_2 vssa1 1.60fF
C789 top_pll_v2_0/div_by_2_0/DFlipFlop_0/CLK vssa1 0.31fF
C790 top_pll_v2_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C791 top_pll_v2_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C792 top_pll_v2_0/div_by_2_0/DFlipFlop_0/nCLK vssa1 1.03fF
C793 top_pll_v2_0/out_div_2 vssa1 -1.30fF
C794 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C795 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C796 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C797 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C798 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C799 top_pll_v2_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C800 top_pll_v2_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C801 top_pll_v2_0/n_out_div_2 vssa1 1.95fF
C802 top_pll_v2_0/div_by_2_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C803 top_pll_v2_0/lf_vc vssa1 -59.89fF
C804 top_pll_v2_0/loop_filter_v2_0/res_loop_filter_2/out vssa1 7.90fF
C805 gpio_noesd[8] vssa1 210.79fF
C806 top_pll_v2_0/loop_filter_v2_0/cap3_loop_filter_0/in vssa1 -12.03fF
C807 top_pll_v2_0/nswitch vssa1 3.73fF
C808 top_pll_v2_0/biasp vssa1 5.44fF
C809 bias_0/iref_1 vssa1 -93.46fF
C810 top_pll_v2_0/vco_vctrl vssa1 -20.08fF
C811 top_pll_v2_0/pswitch vssa1 3.57fF
C812 bias_0/iref_4 vssa1 1.17fF
C813 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219# vssa1 2.60fF
C814 bias_0/iref_3 vssa1 0.64fF
C815 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219# vssa1 2.60fF
C816 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219# vssa1 2.60fF
C817 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219# vssa1 2.60fF
C818 io_analog[5] vssa1 33.29fF
C819 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_0/a_n1731_n1219# vssa1 2.60fF
C820 bias_0/m1_20168_984# vssa1 56.92fF
C821 bias_0/iref_9 vssa1 -1.13fF
C822 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219# vssa1 2.60fF
C823 bias_0/iref_7 vssa1 -1.38fF
C824 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219# vssa1 2.60fF
C825 bias_0/iref_8 vssa1 -1.19fF
C826 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219# vssa1 2.60fF
C827 bias_0/iref_6 vssa1 -1.00fF
C828 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219# vssa1 2.60fF
C829 bias_0/iref_5 vssa1 1.40fF
C830 bias_0/sky130_fd_pr__pfet_01v8_lvt_8P223X_6/a_n1731_n1219# vssa1 2.60fF
C831 top_pll_v1_1/PFD_0/and_pfd_0/a_656_410# vssa1 0.96fF
C832 top_pll_v1_1/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vssa1 0.05fF
C833 top_pll_v1_1/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vssa1 0.05fF
C834 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C835 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_2/B vssa1 1.40fF
C836 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C837 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_3/A vssa1 3.14fF
C838 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C839 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C840 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_2/A vssa1 2.55fF
C841 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C842 top_pll_v1_1/QB vssa1 4.35fF
C843 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C844 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C845 top_pll_v1_1/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C846 top_pll_v1_1/out_div_by_5 vssa1 -0.40fF
C847 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C848 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_2/B vssa1 1.40fF
C849 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C850 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_3/A vssa1 3.14fF
C851 top_pll_v1_1/pfd_reset vssa1 2.17fF
C852 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C853 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C854 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_2/A vssa1 2.55fF
C855 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C856 top_pll_v1_1/QA vssa1 4.22fF
C857 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C858 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C859 top_pll_v1_1/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C860 io_analog[10] vssa1 503.33fF
C861 top_pll_v1_1/pfd_cp_interface_0/inverter_cp_x1_2/in vssa1 1.85fF
C862 top_pll_v1_1/pfd_cp_interface_0/inverter_cp_x1_0/out vssa1 1.77fF
C863 top_pll_v1_1/nUp vssa1 5.39fF
C864 top_pll_v1_1/Up vssa1 1.85fF
C865 top_pll_v1_1/Down vssa1 6.19fF
C866 top_pll_v1_1/nDown vssa1 -3.53fF
C867 top_pll_v1_1/div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vssa1 0.37fF
C868 top_pll_v1_1/div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vssa1 0.38fF
C869 top_pll_v1_1/div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vssa1 0.38fF
C870 top_pll_v1_1/div_by_5_0/DFlipFlop_3/nQ vssa1 0.48fF
C871 top_pll_v1_1/div_5_Q1_shift vssa1 -0.14fF
C872 top_pll_v1_1/div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vssa1 0.57fF
C873 top_pll_v1_1/div_by_5_0/DFlipFlop_3/latch_diff_1/nD vssa1 0.57fF
C874 top_pll_v1_1/div_by_5_0/DFlipFlop_3/latch_diff_1/D vssa1 -1.73fF
C875 top_pll_v1_1/div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vssa1 0.57fF
C876 top_pll_v1_1/div_by_5_0/DFlipFlop_3/latch_diff_0/D vssa1 0.96fF
C877 top_pll_v1_1/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C878 top_pll_v1_1/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C879 top_pll_v1_1/div_by_5_0/DFlipFlop_3/latch_diff_0/nD vssa1 1.14fF
C880 top_pll_v1_1/div_by_5_0/DFlipFlop_2/nQ vssa1 0.48fF
C881 top_pll_v1_1/div_5_Q1 vssa1 4.25fF
C882 top_pll_v1_1/div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vssa1 0.57fF
C883 top_pll_v1_1/div_by_5_0/DFlipFlop_2/latch_diff_1/nD vssa1 0.57fF
C884 top_pll_v1_1/div_by_5_0/DFlipFlop_2/latch_diff_1/D vssa1 -1.73fF
C885 top_pll_v1_1/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vssa1 0.57fF
C886 top_pll_v1_1/div_by_5_0/DFlipFlop_2/latch_diff_0/D vssa1 0.96fF
C887 top_pll_v1_1/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C888 top_pll_v1_1/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C889 top_pll_v1_1/div_by_5_0/DFlipFlop_2/D vssa1 3.13fF
C890 top_pll_v1_1/div_by_5_0/DFlipFlop_2/latch_diff_0/nD vssa1 1.14fF
C891 top_pll_v1_1/div_5_nQ0 vssa1 0.59fF
C892 top_pll_v1_1/div_5_Q0 vssa1 0.01fF
C893 top_pll_v1_1/div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vssa1 0.57fF
C894 top_pll_v1_1/div_by_5_0/DFlipFlop_1/latch_diff_1/nD vssa1 0.57fF
C895 top_pll_v1_1/div_by_5_0/DFlipFlop_1/latch_diff_1/D vssa1 -1.73fF
C896 top_pll_v1_1/div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vssa1 0.57fF
C897 top_pll_v1_1/div_by_5_0/DFlipFlop_1/latch_diff_0/D vssa1 0.96fF
C898 top_pll_v1_1/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C899 top_pll_v1_1/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C900 top_pll_v1_1/div_by_5_0/DFlipFlop_1/D vssa1 3.64fF
C901 top_pll_v1_1/div_by_5_0/DFlipFlop_1/latch_diff_0/nD vssa1 1.14fF
C902 top_pll_v1_1/div_5_nQ2 vssa1 1.24fF
C903 top_pll_v1_1/div_by_5_0/DFlipFlop_0/Q vssa1 -0.94fF
C904 top_pll_v1_1/div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C905 top_pll_v1_1/n_out_by_2 vssa1 -2.75fF
C906 top_pll_v1_1/div_by_5_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C907 top_pll_v1_1/div_by_5_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C908 top_pll_v1_1/div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C909 top_pll_v1_1/out_by_2 vssa1 -5.01fF
C910 top_pll_v1_1/div_by_5_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C911 top_pll_v1_1/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C912 top_pll_v1_1/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C913 top_pll_v1_1/div_by_5_0/DFlipFlop_0/D vssa1 3.96fF
C914 top_pll_v1_1/div_by_5_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C915 top_pll_v1_1/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vssa1 0.08fF
C916 top_pll_v1_1/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vssa1 0.40fF
C917 top_pll_v1_1/out_to_buffer vssa1 1.54fF
C918 top_pll_v1_1/out_to_div vssa1 4.23fF
C919 top_pll_v1_1/out_first_buffer vssa1 2.88fF
C920 top_pll_v1_1/ring_osc_0/csvco_branch_2/in vssa1 1.60fF
C921 top_pll_v1_1/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vssa1 0.16fF
C922 top_pll_v1_1/ring_osc_0/csvco_branch_1/cap_vco_0/t vssa1 7.10fF
C923 top_pll_v1_1/ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vssa1 0.52fF
C924 top_pll_v1_1/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vssa1 0.16fF
C925 top_pll_v1_1/ring_osc_0/csvco_branch_2/cap_vco_0/t vssa1 7.10fF
C926 top_pll_v1_1/ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vssa1 0.52fF
C927 top_pll_v1_1/ring_osc_0/csvco_branch_1/in vssa1 1.58fF
C928 top_pll_v1_1/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vssa1 0.16fF
C929 top_pll_v1_1/vco_out vssa1 1.01fF
C930 top_pll_v1_1/ring_osc_0/csvco_branch_0/cap_vco_0/t vssa1 7.10fF
C931 top_pll_v1_1/ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vssa1 0.52fF
C932 top_pll_v1_1/ring_osc_0/csvco_branch_2/vbp vssa1 0.36fF
C933 io_analog[7] vssa1 24.61fF
C934 top_pll_v1_1/buffer_salida_0/a_3996_n100# vssa1 48.11fF
C935 top_pll_v1_1/buffer_salida_0/a_678_n100# vssa1 13.21fF
C936 top_pll_v1_1/n_out_buffer_div_2 vssa1 1.63fF
C937 top_pll_v1_1/out_buffer_div_2 vssa1 1.60fF
C938 top_pll_v1_1/div_by_2_0/DFlipFlop_0/CLK vssa1 0.31fF
C939 top_pll_v1_1/div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C940 top_pll_v1_1/div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C941 top_pll_v1_1/div_by_2_0/DFlipFlop_0/nCLK vssa1 1.03fF
C942 top_pll_v1_1/out_div_2 vssa1 -1.30fF
C943 top_pll_v1_1/div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C944 top_pll_v1_1/div_by_2_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C945 top_pll_v1_1/div_by_2_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C946 top_pll_v1_1/div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C947 top_pll_v1_1/div_by_2_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C948 top_pll_v1_1/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C949 top_pll_v1_1/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C950 top_pll_v1_1/n_out_div_2 vssa1 1.95fF
C951 top_pll_v1_1/div_by_2_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C952 top_pll_v1_1/nswitch vssa1 3.73fF
C953 top_pll_v1_1/biasp vssa1 5.44fF
C954 bias_0/iref_0 vssa1 -81.35fF
C955 top_pll_v1_1/vco_vctrl vssa1 -18.17fF
C956 top_pll_v1_1/pswitch vssa1 3.57fF
C957 top_pll_v1_1/lf_vc vssa1 -59.89fF
C958 top_pll_v1_1/loop_filter_0/res_loop_filter_2/out vssa1 7.90fF
C959 top_pll_v1_0/PFD_0/and_pfd_0/a_656_410# vssa1 0.96fF
C960 top_pll_v1_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_63_n45# vssa1 0.05fF
C961 top_pll_v1_0/PFD_0/and_pfd_0/sky130_fd_pr__nfet_01v8_ZCYAJJ_0/a_n129_n45# vssa1 0.05fF
C962 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C963 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_2/B vssa1 1.40fF
C964 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C965 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_3/A vssa1 3.14fF
C966 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C967 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C968 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_2/A vssa1 2.55fF
C969 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C970 top_pll_v1_0/QB vssa1 4.35fF
C971 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C972 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C973 top_pll_v1_0/PFD_0/dff_pfd_1/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C974 top_pll_v1_0/out_div_by_5 vssa1 -0.40fF
C975 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C976 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_2/B vssa1 1.40fF
C977 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_3/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C978 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_3/A vssa1 3.14fF
C979 top_pll_v1_0/pfd_reset vssa1 2.17fF
C980 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C981 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_2/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C982 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_2/A vssa1 2.55fF
C983 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C984 top_pll_v1_0/QA vssa1 4.22fF
C985 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_1/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C986 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_63_n90# vssa1 0.03fF
C987 top_pll_v1_0/PFD_0/dff_pfd_0/nor_pfd_0/sky130_fd_pr__pfet_01v8_4F35BC_0/a_n129_n90# vssa1 0.03fF
C988 top_pll_v1_0/pfd_cp_interface_0/inverter_cp_x1_2/in vssa1 1.85fF
C989 top_pll_v1_0/pfd_cp_interface_0/inverter_cp_x1_0/out vssa1 1.77fF
C990 top_pll_v1_0/nUp vssa1 5.39fF
C991 top_pll_v1_0/Up vssa1 1.85fF
C992 top_pll_v1_0/Down vssa1 6.19fF
C993 top_pll_v1_0/nDown vssa1 -3.53fF
C994 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__or2_1_0/a_63_368# vssa1 0.37fF
C995 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__and2_1_1/a_56_136# vssa1 0.38fF
C996 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__and2_1_0/a_56_136# vssa1 0.38fF
C997 top_pll_v1_0/div_by_5_0/DFlipFlop_3/nQ vssa1 0.48fF
C998 top_pll_v1_0/div_5_Q1_shift vssa1 -0.14fF
C999 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_1/m1_657_280# vssa1 0.57fF
C1000 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_1/nD vssa1 0.57fF
C1001 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_1/D vssa1 -1.73fF
C1002 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_0/m1_657_280# vssa1 0.57fF
C1003 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_0/D vssa1 0.96fF
C1004 top_pll_v1_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1005 top_pll_v1_0/div_by_5_0/DFlipFlop_3/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1006 top_pll_v1_0/div_by_5_0/DFlipFlop_3/latch_diff_0/nD vssa1 1.14fF
C1007 top_pll_v1_0/div_by_5_0/DFlipFlop_2/nQ vssa1 0.48fF
C1008 top_pll_v1_0/div_5_Q1 vssa1 4.25fF
C1009 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_1/m1_657_280# vssa1 0.57fF
C1010 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_1/nD vssa1 0.57fF
C1011 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_1/D vssa1 -1.73fF
C1012 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_0/m1_657_280# vssa1 0.57fF
C1013 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_0/D vssa1 0.96fF
C1014 top_pll_v1_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1015 top_pll_v1_0/div_by_5_0/DFlipFlop_2/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1016 top_pll_v1_0/div_by_5_0/DFlipFlop_2/D vssa1 3.13fF
C1017 top_pll_v1_0/div_by_5_0/DFlipFlop_2/latch_diff_0/nD vssa1 1.14fF
C1018 top_pll_v1_0/div_5_nQ0 vssa1 0.59fF
C1019 top_pll_v1_0/div_5_Q0 vssa1 0.01fF
C1020 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_1/m1_657_280# vssa1 0.57fF
C1021 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_1/nD vssa1 0.57fF
C1022 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_1/D vssa1 -1.73fF
C1023 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_0/m1_657_280# vssa1 0.57fF
C1024 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_0/D vssa1 0.96fF
C1025 top_pll_v1_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1026 top_pll_v1_0/div_by_5_0/DFlipFlop_1/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1027 top_pll_v1_0/div_by_5_0/DFlipFlop_1/D vssa1 3.64fF
C1028 top_pll_v1_0/div_by_5_0/DFlipFlop_1/latch_diff_0/nD vssa1 1.14fF
C1029 top_pll_v1_0/div_5_nQ2 vssa1 1.24fF
C1030 top_pll_v1_0/div_by_5_0/DFlipFlop_0/Q vssa1 -0.94fF
C1031 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C1032 top_pll_v1_0/n_out_by_2 vssa1 -2.75fF
C1033 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C1034 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C1035 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C1036 top_pll_v1_0/out_by_2 vssa1 -5.01fF
C1037 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C1038 top_pll_v1_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1039 top_pll_v1_0/div_by_5_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1040 top_pll_v1_0/div_by_5_0/DFlipFlop_0/D vssa1 3.96fF
C1041 top_pll_v1_0/div_by_5_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C1042 vdda1 vssa1 6838.97fF
C1043 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_355_368# vssa1 0.08fF
C1044 top_pll_v1_0/div_by_5_0/sky130_fd_sc_hs__xor2_1_0/a_194_125# vssa1 0.40fF
C1045 top_pll_v1_0/out_to_buffer vssa1 1.54fF
C1046 top_pll_v1_0/out_to_div vssa1 4.23fF
C1047 top_pll_v1_0/out_first_buffer vssa1 2.88fF
C1048 top_pll_v1_0/ring_osc_0/csvco_branch_2/in vssa1 1.60fF
C1049 top_pll_v1_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vdd vssa1 0.16fF
C1050 top_pll_v1_0/ring_osc_0/csvco_branch_1/cap_vco_0/t vssa1 7.10fF
C1051 top_pll_v1_0/ring_osc_0/csvco_branch_1/inverter_csvco_0/vss vssa1 0.52fF
C1052 top_pll_v1_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vdd vssa1 0.16fF
C1053 top_pll_v1_0/ring_osc_0/csvco_branch_2/cap_vco_0/t vssa1 7.10fF
C1054 top_pll_v1_0/ring_osc_0/csvco_branch_2/inverter_csvco_0/vss vssa1 0.52fF
C1055 top_pll_v1_0/ring_osc_0/csvco_branch_1/in vssa1 1.58fF
C1056 top_pll_v1_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vdd vssa1 0.16fF
C1057 top_pll_v1_0/vco_out vssa1 1.01fF
C1058 gpio_noesd[7] vssa1 272.21fF
C1059 top_pll_v1_0/ring_osc_0/csvco_branch_0/cap_vco_0/t vssa1 7.10fF
C1060 top_pll_v1_0/ring_osc_0/csvco_branch_0/inverter_csvco_0/vss vssa1 0.52fF
C1061 top_pll_v1_0/ring_osc_0/csvco_branch_2/vbp vssa1 0.36fF
C1062 io_analog[9] vssa1 7.89fF
C1063 top_pll_v1_0/buffer_salida_0/a_3996_n100# vssa1 48.23fF
C1064 top_pll_v1_0/buffer_salida_0/a_678_n100# vssa1 13.21fF
C1065 top_pll_v1_0/n_out_buffer_div_2 vssa1 1.63fF
C1066 top_pll_v1_0/out_buffer_div_2 vssa1 1.60fF
C1067 top_pll_v1_0/div_by_2_0/DFlipFlop_0/CLK vssa1 0.31fF
C1068 top_pll_v1_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1069 top_pll_v1_0/div_by_2_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1070 top_pll_v1_0/div_by_2_0/DFlipFlop_0/nCLK vssa1 1.03fF
C1071 top_pll_v1_0/out_div_2 vssa1 -1.30fF
C1072 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_1/m1_657_280# vssa1 0.57fF
C1073 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_1/nD vssa1 0.57fF
C1074 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_1/D vssa1 -1.73fF
C1075 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_0/m1_657_280# vssa1 0.57fF
C1076 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_0/D vssa1 0.96fF
C1077 top_pll_v1_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_2/in vssa1 1.86fF
C1078 top_pll_v1_0/div_by_2_0/DFlipFlop_0/clock_inverter_0/inverter_cp_x1_0/out vssa1 1.76fF
C1079 top_pll_v1_0/n_out_div_2 vssa1 1.95fF
C1080 top_pll_v1_0/div_by_2_0/DFlipFlop_0/latch_diff_0/nD vssa1 1.14fF
C1081 top_pll_v1_0/nswitch vssa1 3.73fF
C1082 top_pll_v1_0/biasp vssa1 5.44fF
C1083 bias_0/iref_2 vssa1 -186.53fF
C1084 top_pll_v1_0/vco_vctrl vssa1 -18.17fF
C1085 top_pll_v1_0/pswitch vssa1 3.57fF
C1086 top_pll_v1_0/lf_vc vssa1 -59.89fF
C1087 top_pll_v1_0/loop_filter_0/res_loop_filter_2/out vssa1 7.90fF
.ends

