**.subckt tb_prescaler_23
VSS vss GND {vss} 
VDD vdd vss {vdd} 
Vref CLK vss PULSE(0 {vin} 0 1p 1p {Tref/2} {Tref}) DC {vin} AC 0 
C2 clk_23 vss 10f m=1
x2 nclk_2 vss CLK vdd clk_2 net1 net2 net3 net4 div_by_2
x1 vdd clk_23 clk_2 nclk_2 vss MC net6 net5 net7 net8 prescaler_23
VMC MC vss PULSE(0 {vin} 0 1p 1p 400n 800n) DC {vin} AC 0 
**** begin user architecture code



* Parameters
.param kp = 1.0
.param vdd = kp*1.8
.param vss = 0.0
.param vin = vdd
.param fref = 1e9
.param Tref = 1/fref
.param C = 1f
.param iref=100u

.options TEMP = 100.0
.options RSHUNT = 1e20

* Models
.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib SS

* Data to save
.save all
.ic v(CLK) = 0.0
.ic v(MC) = 0.0
.ic v(clk_2) = 0.0
.ic v(nclk_2) = 0.0
.ic v(clk_23) = 0.0

* Simulation
.control
	tran 0.01ns 800ns
	write tb_div_by_5_tran.raw
	plot v(clk_23) v(clk) v(clk_2) v(clk_23)+3 v(clk_2)+6 v(clk)+9

.endc



**** end user architecture code
**.ends

* expanding   symbol:  div_by_2/sch/div_by_2.sym # of pins=9
* sym_path: /home/dhernando/sky130-mpw2-fulgor/div_by_2/sch/div_by_2.sym
* sch_path: /home/dhernando/sky130-mpw2-fulgor/div_by_2/sch/div_by_2.sch
.subckt div_by_2  nCLK_2 vss CLK vdd CLK_2 out_div nout_div o1 o2
*.ipin CLK
*.opin CLK_2
*.iopin vss
*.iopin vdd
*.opin nCLK_2
*.iopin nout_div
*.iopin o2
*.iopin o1
*.iopin out_div
x1 vdd out_div nout_div vss nout_div CLK_d nCLK_d DFlipFlop
x2 vdd CLK_d CLK nCLK_d vss clock_inverter
x3 vdd o1 out_div vss inverter_min_x2
x4 vdd CLK_2 o1 vss inverter_min_x4
x5 vdd o2 nout_div vss inverter_min_x2
x6 vdd nCLK_2 o2 vss inverter_min_x4
.ends


* expanding   symbol:  prescaler_23/sch/prescaler_23.sym # of pins=10
* sym_path: /home/dhernando/sky130-mpw2-fulgor/prescaler_23/sch/prescaler_23.sym
* sch_path: /home/dhernando/sky130-mpw2-fulgor/prescaler_23/sch/prescaler_23.sch
.subckt prescaler_23  vdd CLK_23 CLK nCLK vss MC Q1 nCLK_23 Q2 Q2_d
*.iopin vdd
*.ipin CLK
*.ipin nCLK
*.ipin MC
*.iopin vss
*.opin CLK_23
*.iopin nCLK_23
*.iopin Q1
*.iopin Q2
*.iopin Q2_d
x3 nCLK_23 1 vss vss vdd vdd 2 sky130_fd_sc_hs__and2_1
x4 Q1 MC vss vss vdd vdd 1 sky130_fd_sc_hs__or2_1
x6 3 nCLK_23 MC vss vss vdd vdd CLK_23 sky130_fd_sc_hs__mux2_1
x7 Q2 Q2_d vss vss vdd vdd 3 sky130_fd_sc_hs__or2_1
x1 vdd Q1 net1 vss nCLK_23 CLK nCLK DFlipFlop
x2 vdd Q2 nCLK_23 vss 2 CLK nCLK DFlipFlop
x5 vdd Q2_d net2 vss Q2 nCLK CLK DFlipFlop
.ends


* expanding   symbol:  DFlipFlop/sch/DFlipFlop.sym # of pins=7
* sym_path: /home/dhernando/sky130-mpw2-fulgor/DFlipFlop/sch/DFlipFlop.sym
* sch_path: /home/dhernando/sky130-mpw2-fulgor/DFlipFlop/sch/DFlipFlop.sch
.subckt DFlipFlop  vdd Q nQ vss D CLK nCLK
*.iopin vdd
*.iopin vss
*.opin Q
*.opin nQ
*.ipin D
*.ipin CLK
*.ipin nCLK
x1 vdd D_d D nD_d vss clock_inverter
x2 vdd nA A D_d nD_d CLK vss latch_diff
x3 vdd nQ Q A nA nCLK vss latch_diff
.ends


* expanding   symbol:  clock_inverter/sch/clock_inverter.sym # of pins=5
* sym_path: /home/dhernando/sky130-mpw2-fulgor/clock_inverter/sch/clock_inverter.sym
* sch_path: /home/dhernando/sky130-mpw2-fulgor/clock_inverter/sch/clock_inverter.sch
.subckt clock_inverter  vdd CLK_d CLK nCLK_d vss
*.ipin CLK
*.iopin vdd
*.iopin vss
*.opin nCLK_d
*.opin CLK_d
x5 vdd nCLK_d net1 vss trans_gate
x1 vdd CLK_d net2 vss inverter_cp_x1
x2 vdd net2 CLK vss inverter_cp_x1
x3 vdd net1 CLK vss inverter_cp_x1
.ends


* expanding   symbol:  inverter_min_x2/sch/inverter_min_x2.sym # of pins=4
* sym_path: /home/dhernando/sky130-mpw2-fulgor/inverter_min_x2/sch/inverter_min_x2.sym
* sch_path: /home/dhernando/sky130-mpw2-fulgor/inverter_min_x2/sch/inverter_min_x2.sch
.subckt inverter_min_x2  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:  inverter_min_x4/sch/inverter_min_x4.sym # of pins=4
* sym_path: /home/dhernando/sky130-mpw2-fulgor/inverter_min_x4/sch/inverter_min_x4.sym
* sch_path: /home/dhernando/sky130-mpw2-fulgor/inverter_min_x4/sch/inverter_min_x4.sch
.subckt inverter_min_x4  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
.ends


* expanding   symbol:  latch_diff/sch/latch_diff.sym # of pins=7
* sym_path: /home/dhernando/sky130-mpw2-fulgor/latch_diff/sch/latch_diff.sym
* sch_path: /home/dhernando/sky130-mpw2-fulgor/latch_diff/sch/latch_diff.sch
.subckt latch_diff  vdd nQ Q D nD CLK vss
*.iopin vdd
*.iopin vss
*.ipin D
*.opin nQ
*.ipin CLK
*.ipin nD
*.opin Q
XM3 net1 CLK vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM4 nQ Q vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM5 Q nQ vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM1 nQ D net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 Q nD net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.95 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:  trans_gate/sch/trans_gate.sym # of pins=4
* sym_path: /home/dhernando/sky130-mpw2-fulgor/trans_gate/sch/trans_gate.sym
* sch_path: /home/dhernando/sky130-mpw2-fulgor/trans_gate/sch/trans_gate.sch
.subckt trans_gate  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out vss in vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM1 out vdd in vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
.ends


* expanding   symbol:  inverter_cp_x1/sch/inverter_cp_x1.sym # of pins=4
* sym_path: /home/dhernando/sky130-mpw2-fulgor/inverter_cp_x1/sch/inverter_cp_x1.sym
* sch_path: /home/dhernando/sky130-mpw2-fulgor/inverter_cp_x1/sch/inverter_cp_x1.sch
.subckt inverter_cp_x1  vdd out in vss
*.iopin vss
*.ipin in
*.opin out
*.iopin vdd
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
.ends

.GLOBAL GND
**** begin user architecture code
.include ~/skywater/skywater-pdk/libraries/sky130_fd_sc_hs/latest/cells/and2/sky130_fd_sc_hs__and2_1.spice
.include ~/skywater/skywater-pdk/libraries/sky130_fd_sc_hs/latest/cells/or2/sky130_fd_sc_hs__or2_1.spice
.include ~/skywater/skywater-pdk/libraries/sky130_fd_sc_hs/latest/cells/mux2/sky130_fd_sc_hs__mux2_1.spice

**** end user architecture code
** flattened .save nodes
.end
