magic
tech sky130A
magscale 1 2
timestamp 1624022177
<< pwell >>
rect -16462 -24206 34360 5780
<< psubdiff >>
rect -16450 4360 -14850 4384
rect -16450 -21664 -14850 -21640
rect 32749 4360 34349 4384
rect -16450 -22594 -14851 -21664
rect 32749 -22593 34349 -21640
rect 32749 -22594 34348 -22593
rect -16450 -24194 -11039 -22594
rect 28961 -24194 34348 -22594
<< psubdiffcont >>
rect -16450 -21640 -14850 4360
rect 32749 -21640 34349 4360
rect -11039 -24194 28961 -22594
<< locali >>
rect -16450 4360 -14850 4376
rect 32749 4360 34349 4376
rect -14851 -21656 -14850 -21640
rect 34348 -21656 34349 -21640
<< viali >>
rect -16450 -21640 -14850 4360
rect 135 -119 4328 -40
rect -16450 -22594 -14851 -21640
rect 32749 -21640 34349 4360
rect 32749 -22594 34348 -21640
rect -16450 -24194 -11039 -22594
rect -11039 -24194 28961 -22594
rect 28961 -24194 34348 -22594
<< metal1 >>
rect -370 5080 -360 5680
rect 640 5614 650 5680
rect 2456 5614 2466 5680
rect 640 5182 1312 5614
rect 1560 5182 2466 5614
rect 640 5080 650 5182
rect 2456 5080 2466 5182
rect 3866 5614 3876 5680
rect 3866 5182 4100 5614
rect 3866 5080 3876 5182
rect -16456 4360 -14844 4372
rect -16456 -21634 -16450 4360
rect -16462 -24194 -16450 -21634
rect -14850 -21634 -14844 4360
rect 32743 4360 34355 4372
rect 166 166 3245 598
rect 40 -40 4361 83
rect 40 -119 135 -40
rect 4328 -119 4361 -40
rect 40 -213 4361 -119
rect 1312 -1221 2954 -213
rect 1312 -1273 2955 -1221
rect 1313 -2326 2955 -1273
rect -14850 -21640 -14839 -21634
rect -14851 -22588 -14839 -21640
rect 1313 -22588 2954 -2326
rect 32743 -22588 32749 4360
rect 34349 -21640 34355 4360
rect -14851 -22594 32749 -22588
rect 34348 -21652 34355 -21640
rect 34348 -22588 34354 -21652
rect 34348 -24194 34360 -22588
rect -16462 -24200 34360 -24194
rect 32743 -24206 34354 -24200
<< via1 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -10029 -23953 -4329 -22753
rect 9433 -24034 31413 -22834
<< metal2 >>
rect -360 5680 640 5690
rect -360 5070 640 5080
rect 2466 5680 3866 5690
rect 2466 5070 3866 5080
rect -10029 -22753 -4329 -22743
rect -10029 -23963 -4329 -23953
rect 9433 -22834 31413 -22824
rect 9433 -24044 31413 -24034
<< via2 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
rect -10029 -23953 -4329 -22753
rect 9433 -24034 31413 -22834
<< metal3 >>
rect -370 5680 650 5685
rect -370 5080 -360 5680
rect 640 5080 650 5680
rect -370 5075 650 5080
rect 2456 5680 3876 5685
rect 2456 5080 2466 5680
rect 3866 5080 3876 5680
rect 2456 5075 3876 5080
rect -10059 -22753 -4267 -9184
rect 4852 -21602 9433 4898
rect 10833 -21602 14842 4898
rect 16242 -21602 20055 4898
rect 21455 -21602 25394 4898
rect 26794 -21602 31427 4898
rect -10059 -23008 -10029 -22753
rect -10039 -23953 -10029 -23008
rect -4329 -23008 -4267 -22753
rect 30027 -22829 31427 -21602
rect -4329 -23136 -4295 -23008
rect -4329 -23953 -4319 -23136
rect -10039 -23958 -4319 -23953
rect 9423 -24034 9433 -22829
rect 10833 -22834 14842 -22829
rect 16242 -22834 20055 -22829
rect 21455 -22834 25394 -22829
rect 26794 -22834 31427 -22829
rect 31413 -23602 31427 -22834
rect 31413 -24034 31423 -23602
rect 9423 -24039 31423 -24034
rect 25394 -24061 26794 -24039
<< via3 >>
rect -360 5080 640 5680
rect 2466 5080 3866 5680
<< metal4 >>
rect -10754 5680 740 5780
rect -10754 5080 -360 5680
rect 640 5080 740 5680
rect -10754 4980 740 5080
rect 2066 5680 28119 5780
rect 2066 5080 2466 5680
rect 3866 5080 28119 5680
rect 2066 4980 28119 5080
use cap2_loop_filter  cap2_loop_filter_0
timestamp 1624021628
transform 1 0 -4885 0 1 288
box -8638 -9892 4299 5492
use cap1_loop_filter  cap1_loop_filter_0
timestamp 1624018159
transform 1 0 47404 0 1 20622
box -42552 -43690 -15977 -14842
use res_loop_filter  res_loop_filter_0
timestamp 1624015667
transform 1 0 0 0 1 0
box 0 0 1478 5780
use res_loop_filter  res_loop_filter_1
timestamp 1624015667
transform 1 0 1478 0 1 0
box 0 0 1478 5780
use res_loop_filter  res_loop_filter_2
timestamp 1624015667
transform 1 0 2956 0 1 0
box 0 0 1478 5780
<< labels >>
rlabel pwell 1313 -22594 2954 -168 1 vss
rlabel metal4 -10754 4980 -360 5780 1 in
rlabel metal4 3866 4980 28119 5780 1 vc_pex
<< end >>
