magic
tech sky130A
magscale 1 2
timestamp 1624113259
<< nwell >>
rect 291 1100 1333 1369
<< pwell >>
rect -576 -643 2878 -503
<< psubdiff >>
rect -468 -652 -444 -595
rect 2746 -652 2770 -595
<< nsubdiff >>
rect 387 1217 423 1319
rect 685 1217 843 1319
rect 1201 1217 1231 1319
<< psubdiffcont >>
rect -444 -652 2746 -595
<< nsubdiffcont >>
rect 423 1217 685 1319
rect 843 1217 1201 1319
<< viali >>
rect 387 1217 423 1319
rect 423 1217 685 1319
rect 685 1217 843 1319
rect 843 1217 1201 1319
rect 1201 1217 1231 1319
rect 327 1129 1297 1163
rect -540 -595 2842 -503
rect -540 -652 -444 -595
rect -444 -652 2746 -595
rect 2746 -652 2842 -595
<< metal1 >>
rect 281 1359 1343 1369
rect 281 1122 291 1359
rect 1333 1122 1343 1359
rect 511 801 521 980
rect 587 801 597 980
rect 835 801 845 980
rect 911 801 921 980
rect 951 977 997 1122
rect 1027 801 1037 980
rect 1103 801 1113 980
rect 1143 978 1189 1122
rect 435 749 481 791
rect 627 749 673 791
rect 435 739 673 749
rect 435 682 473 739
rect 635 682 673 739
rect 435 670 673 682
rect 1080 674 1090 739
rect 1185 674 1195 739
rect -432 389 2692 525
rect -432 350 -386 389
rect -240 351 -194 389
rect -48 351 -2 389
rect 128 383 2690 389
rect 144 351 190 383
rect -356 151 -346 351
rect -280 151 -270 351
rect -164 151 -154 351
rect -88 151 -78 351
rect 28 151 38 351
rect 104 151 114 351
rect 352 259 362 351
rect 428 259 438 351
rect 544 259 554 351
rect 620 259 630 351
rect 868 259 878 351
rect 944 259 954 351
rect 1060 259 1070 351
rect 1136 259 1146 351
rect 1288 259 1298 351
rect 1364 259 1374 351
rect 1480 259 1490 351
rect 1556 259 1566 351
rect 1672 259 1682 351
rect 1748 259 1758 351
rect 1900 259 1910 351
rect 1976 259 1986 351
rect 2092 259 2102 351
rect 2168 259 2178 351
rect 2284 259 2294 351
rect 2360 259 2370 351
rect 2476 259 2486 351
rect 2552 259 2562 351
rect 2668 259 2678 351
rect 2744 259 2754 351
rect 448 125 458 217
rect 524 125 534 217
rect 640 125 650 217
rect 716 125 726 217
rect 964 125 974 217
rect 1040 125 1050 217
rect 1384 125 1394 217
rect 1460 125 1470 217
rect 1576 125 1586 217
rect 1652 125 1662 217
rect 1996 125 2006 217
rect 2072 125 2082 217
rect 2188 125 2198 217
rect 2264 125 2274 217
rect 2380 125 2390 217
rect 2456 125 2466 217
rect 2572 125 2582 217
rect 2648 125 2658 217
rect 1185 -19 1195 72
rect 1267 -19 1277 72
rect 1809 68 1863 71
rect 239 -85 249 -70
rect 146 -131 249 -85
rect 239 -147 249 -131
rect 315 -85 325 -70
rect 1198 -81 1252 -19
rect 1789 -23 1799 68
rect 1871 -23 1881 68
rect 2788 -16 2798 75
rect 2870 -16 2880 75
rect 1809 -80 1863 -23
rect 2806 -80 2860 -16
rect 315 -131 426 -85
rect 315 -147 325 -131
rect 1067 -135 1252 -81
rect 1682 -134 1863 -80
rect 2658 -134 2860 -80
rect -356 -363 -346 -163
rect -280 -363 -270 -163
rect -164 -363 -154 -163
rect -88 -363 -78 -163
rect 28 -363 38 -163
rect 104 -363 114 -163
rect -432 -497 -386 -363
rect -240 -497 -194 -363
rect -48 -497 -2 -363
rect 144 -497 190 -363
rect 372 -497 418 -357
rect 448 -363 458 -163
rect 524 -363 534 -163
rect 564 -497 610 -357
rect 640 -363 650 -163
rect 716 -363 726 -163
rect 888 -497 934 -359
rect 964 -363 974 -163
rect 1040 -363 1050 -163
rect 1080 -497 1126 -359
rect 1308 -497 1354 -357
rect 1384 -363 1394 -163
rect 1460 -363 1470 -163
rect 1500 -497 1546 -358
rect 1576 -363 1586 -163
rect 1652 -363 1662 -163
rect 1692 -497 1738 -358
rect 1920 -497 1966 -360
rect 1996 -363 2006 -163
rect 2072 -363 2082 -163
rect 2112 -497 2158 -358
rect 2188 -363 2198 -163
rect 2264 -363 2274 -163
rect 2304 -497 2350 -356
rect 2380 -363 2390 -163
rect 2456 -363 2466 -163
rect 2496 -497 2542 -358
rect 2572 -363 2582 -163
rect 2648 -363 2658 -163
rect 2688 -497 2734 -355
rect -586 -676 -576 -497
rect 2878 -676 2888 -497
<< via1 >>
rect 291 1319 1333 1359
rect 291 1217 387 1319
rect 387 1217 1231 1319
rect 1231 1217 1333 1319
rect 291 1163 1333 1217
rect 291 1129 327 1163
rect 327 1129 1297 1163
rect 1297 1129 1333 1163
rect 291 1122 1333 1129
rect 521 801 587 980
rect 845 801 911 980
rect 1037 801 1103 980
rect 473 682 635 739
rect 1090 674 1185 739
rect -346 151 -280 351
rect -154 151 -88 351
rect 38 151 104 351
rect 362 259 428 351
rect 554 259 620 351
rect 878 259 944 351
rect 1070 259 1136 351
rect 1298 259 1364 351
rect 1490 259 1556 351
rect 1682 259 1748 351
rect 1910 259 1976 351
rect 2102 259 2168 351
rect 2294 259 2360 351
rect 2486 259 2552 351
rect 2678 259 2744 351
rect 458 125 524 217
rect 650 125 716 217
rect 974 125 1040 217
rect 1394 125 1460 217
rect 1586 125 1652 217
rect 2006 125 2072 217
rect 2198 125 2264 217
rect 2390 125 2456 217
rect 2582 125 2648 217
rect 1195 -19 1267 72
rect 249 -147 315 -70
rect 1799 -23 1871 68
rect 2798 -16 2870 75
rect -346 -363 -280 -163
rect -154 -363 -88 -163
rect 38 -363 104 -163
rect 458 -363 524 -163
rect 650 -363 716 -163
rect 974 -363 1040 -163
rect 1394 -363 1460 -163
rect 1586 -363 1652 -163
rect 2006 -363 2072 -163
rect 2198 -363 2264 -163
rect 2390 -363 2456 -163
rect 2582 -363 2648 -163
rect -576 -503 2878 -497
rect -576 -652 -540 -503
rect -540 -652 2842 -503
rect 2842 -652 2878 -503
rect -576 -676 2878 -652
<< metal2 >>
rect 249 1359 1333 1369
rect 249 1122 291 1359
rect 249 1112 1333 1122
rect -346 351 -280 361
rect -154 351 -88 361
rect -280 167 -154 340
rect -346 -163 -280 151
rect 38 351 104 361
rect -88 167 38 340
rect -154 -163 -88 151
rect -280 -354 -154 -181
rect -346 -373 -280 -363
rect 38 -163 104 151
rect 249 -70 315 1112
rect 521 980 587 990
rect 845 980 911 990
rect 1037 980 1103 990
rect 587 801 845 980
rect 911 801 1037 980
rect 521 791 587 801
rect 845 791 911 801
rect 1037 791 1103 801
rect 473 739 795 749
rect 635 682 795 739
rect 473 660 795 682
rect 1090 739 1185 749
rect 1090 664 1185 674
rect 362 351 428 361
rect 554 351 620 361
rect 682 351 795 660
rect 878 351 944 361
rect 1070 351 1136 361
rect 1298 351 1364 361
rect 1490 351 1556 361
rect 1682 351 1748 361
rect 1910 351 1976 361
rect 2102 351 2168 361
rect 2294 351 2360 361
rect 2486 351 2552 361
rect 2678 351 2744 361
rect 428 259 554 351
rect 620 259 878 351
rect 944 259 1070 351
rect 1136 259 1298 351
rect 1364 259 1490 351
rect 1556 259 1682 351
rect 1748 259 1910 351
rect 1976 259 2102 351
rect 2168 259 2294 351
rect 2360 259 2486 351
rect 2552 259 2678 351
rect 362 249 428 259
rect 554 249 620 259
rect 878 249 944 259
rect 1070 249 1136 259
rect 1298 249 1364 259
rect 1490 249 1556 259
rect 1682 249 1748 259
rect 1910 249 1976 259
rect 2102 249 2168 259
rect 2294 249 2360 259
rect 2486 249 2552 259
rect 2678 249 2744 259
rect 249 -157 315 -147
rect 458 217 524 227
rect 650 217 716 227
rect 524 154 650 199
rect -88 -354 38 -181
rect -154 -373 -88 -363
rect 38 -373 104 -363
rect 458 -163 524 125
rect 650 -163 716 125
rect 524 -363 650 -163
rect 458 -373 524 -363
rect 650 -373 716 -363
rect 974 217 1040 227
rect 974 -163 1040 125
rect 1394 217 1460 227
rect 1195 72 1267 82
rect 1195 -29 1267 -19
rect 974 -373 1040 -363
rect 1394 -163 1460 125
rect 1586 217 1652 227
rect 1586 -163 1652 125
rect 2006 217 2072 227
rect 1799 68 1871 78
rect 1799 -33 1871 -23
rect 1460 -363 1586 -163
rect 1394 -373 1460 -363
rect 1586 -373 1652 -363
rect 2006 -163 2072 125
rect 2198 217 2264 227
rect 2198 -163 2264 125
rect 2390 217 2456 227
rect 2390 -163 2456 125
rect 2582 217 2648 227
rect 2582 -163 2648 125
rect 2798 75 2870 85
rect 2798 -26 2870 -16
rect 2072 -363 2198 -163
rect 2264 -363 2390 -163
rect 2456 -363 2582 -163
rect 2006 -373 2072 -363
rect 2198 -373 2264 -363
rect 2390 -373 2456 -363
rect 2582 -373 2648 -363
rect -576 -497 2878 -487
rect -576 -686 2878 -676
<< via2 >>
rect 1090 674 1185 739
rect 1195 -19 1267 72
rect 1799 -23 1871 68
rect 2798 -16 2870 75
rect 1168 -626 1263 -561
<< metal3 >>
rect 1024 739 1195 744
rect 1024 674 1090 739
rect 1185 674 1195 739
rect 1024 669 1195 674
rect 1024 -556 1114 669
rect 1185 72 1279 82
rect 1185 -19 1195 72
rect 1267 -19 1279 72
rect 1185 -24 1279 -19
rect 1789 68 1883 78
rect 1789 -23 1799 68
rect 1871 -23 1883 68
rect 2788 75 2882 85
rect 2788 -16 2798 75
rect 2870 -16 2882 75
rect 2788 -21 2882 -16
rect 1789 -28 1883 -23
rect 1024 -561 1273 -556
rect 1024 -626 1168 -561
rect 1263 -626 1273 -561
rect 1024 -631 1273 -626
use sky130_fd_pr__nfet_01v8_lvt_9B2JY7  sky130_fd_pr__nfet_01v8_lvt_9B2JY7_0
timestamp 1624020979
transform 1 0 -121 0 1 251
box -455 -310 455 310
use sky130_fd_pr__nfet_01v8_lvt_9B2JY7  sky130_fd_pr__nfet_01v8_lvt_9B2JY7_1
timestamp 1624020979
transform 1 0 -121 0 1 -263
box -455 -310 455 310
use sky130_fd_pr__nfet_01v8_lvt_72JNYZ  sky130_fd_pr__nfet_01v8_lvt_72JNYZ_1
timestamp 1624032293
transform 1 0 539 0 1 -263
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_lvt_72JNYZ  sky130_fd_pr__nfet_01v8_lvt_72JNYZ_0
timestamp 1624032293
transform 1 0 539 0 1 251
box -311 -310 311 310
use sky130_fd_pr__nfet_01v8_lvt_B2JNY3  sky130_fd_pr__nfet_01v8_lvt_B2JNY3_1
timestamp 1623958660
transform 1 0 1523 0 1 -263
box -359 -310 359 310
use sky130_fd_pr__nfet_01v8_lvt_B2JNY3  sky130_fd_pr__nfet_01v8_lvt_B2JNY3_0
timestamp 1623958660
transform 1 0 1523 0 1 251
box -359 -310 359 310
use sky130_fd_pr__nfet_01v8_lvt_MVT43V  sky130_fd_pr__nfet_01v8_lvt_MVT43V_1
timestamp 1623958102
transform 1 0 1007 0 1 -263
box -263 -310 263 310
use sky130_fd_pr__nfet_01v8_lvt_MVT43V  sky130_fd_pr__nfet_01v8_lvt_MVT43V_0
timestamp 1623958102
transform 1 0 1007 0 1 251
box -263 -310 263 310
use sky130_fd_pr__nfet_01v8_lvt_NMSMYT  sky130_fd_pr__nfet_01v8_lvt_NMSMYT_1
timestamp 1623958459
transform 1 0 2327 0 1 -263
box -551 -310 551 310
use sky130_fd_pr__nfet_01v8_lvt_NMSMYT  sky130_fd_pr__nfet_01v8_lvt_NMSMYT_0
timestamp 1623958459
transform 1 0 2327 0 1 251
box -551 -310 551 310
use sky130_fd_pr__pfet_01v8_XACJHL  sky130_fd_pr__pfet_01v8_XACJHL_0
timestamp 1624020979
transform -1 0 554 0 1 880
box -263 -319 263 319
use sky130_fd_pr__pfet_01v8_XAYTAL  sky130_fd_pr__pfet_01v8_XAYTAL_0
timestamp 1623959550
transform -1 0 1022 0 1 880
box -311 -319 311 319
<< labels >>
rlabel via1 1258 1198 1292 1233 1 avdd1p8
rlabel via1 -540 -584 -506 -549 1 avss1p8
rlabel metal1 168 388 202 423 1 iref
rlabel metal2 739 441 773 476 1 vctrl
rlabel metal3 1215 9 1249 44 1 reg0
rlabel metal3 1819 10 1853 45 1 reg1
rlabel metal3 2809 13 2843 48 1 reg2
<< end >>
