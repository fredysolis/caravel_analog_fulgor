magic
tech sky130A
magscale 1 2
timestamp 1623774805
<< nwell >>
rect -1367 -369 1367 369
<< pmos >>
rect -1167 -150 -1137 150
rect -1071 -150 -1041 150
rect -975 -150 -945 150
rect -879 -150 -849 150
rect -783 -150 -753 150
rect -687 -150 -657 150
rect -591 -150 -561 150
rect -495 -150 -465 150
rect -399 -150 -369 150
rect -303 -150 -273 150
rect -207 -150 -177 150
rect -111 -150 -81 150
rect -15 -150 15 150
rect 81 -150 111 150
rect 177 -150 207 150
rect 273 -150 303 150
rect 369 -150 399 150
rect 465 -150 495 150
rect 561 -150 591 150
rect 657 -150 687 150
rect 753 -150 783 150
rect 849 -150 879 150
rect 945 -150 975 150
rect 1041 -150 1071 150
rect 1137 -150 1167 150
<< pdiff >>
rect -1229 138 -1167 150
rect -1229 -138 -1217 138
rect -1183 -138 -1167 138
rect -1229 -150 -1167 -138
rect -1137 138 -1071 150
rect -1137 -138 -1121 138
rect -1087 -138 -1071 138
rect -1137 -150 -1071 -138
rect -1041 138 -975 150
rect -1041 -138 -1025 138
rect -991 -138 -975 138
rect -1041 -150 -975 -138
rect -945 138 -879 150
rect -945 -138 -929 138
rect -895 -138 -879 138
rect -945 -150 -879 -138
rect -849 138 -783 150
rect -849 -138 -833 138
rect -799 -138 -783 138
rect -849 -150 -783 -138
rect -753 138 -687 150
rect -753 -138 -737 138
rect -703 -138 -687 138
rect -753 -150 -687 -138
rect -657 138 -591 150
rect -657 -138 -641 138
rect -607 -138 -591 138
rect -657 -150 -591 -138
rect -561 138 -495 150
rect -561 -138 -545 138
rect -511 -138 -495 138
rect -561 -150 -495 -138
rect -465 138 -399 150
rect -465 -138 -449 138
rect -415 -138 -399 138
rect -465 -150 -399 -138
rect -369 138 -303 150
rect -369 -138 -353 138
rect -319 -138 -303 138
rect -369 -150 -303 -138
rect -273 138 -207 150
rect -273 -138 -257 138
rect -223 -138 -207 138
rect -273 -150 -207 -138
rect -177 138 -111 150
rect -177 -138 -161 138
rect -127 -138 -111 138
rect -177 -150 -111 -138
rect -81 138 -15 150
rect -81 -138 -65 138
rect -31 -138 -15 138
rect -81 -150 -15 -138
rect 15 138 81 150
rect 15 -138 31 138
rect 65 -138 81 138
rect 15 -150 81 -138
rect 111 138 177 150
rect 111 -138 127 138
rect 161 -138 177 138
rect 111 -150 177 -138
rect 207 138 273 150
rect 207 -138 223 138
rect 257 -138 273 138
rect 207 -150 273 -138
rect 303 138 369 150
rect 303 -138 319 138
rect 353 -138 369 138
rect 303 -150 369 -138
rect 399 138 465 150
rect 399 -138 415 138
rect 449 -138 465 138
rect 399 -150 465 -138
rect 495 138 561 150
rect 495 -138 511 138
rect 545 -138 561 138
rect 495 -150 561 -138
rect 591 138 657 150
rect 591 -138 607 138
rect 641 -138 657 138
rect 591 -150 657 -138
rect 687 138 753 150
rect 687 -138 703 138
rect 737 -138 753 138
rect 687 -150 753 -138
rect 783 138 849 150
rect 783 -138 799 138
rect 833 -138 849 138
rect 783 -150 849 -138
rect 879 138 945 150
rect 879 -138 895 138
rect 929 -138 945 138
rect 879 -150 945 -138
rect 975 138 1041 150
rect 975 -138 991 138
rect 1025 -138 1041 138
rect 975 -150 1041 -138
rect 1071 138 1137 150
rect 1071 -138 1087 138
rect 1121 -138 1137 138
rect 1071 -150 1137 -138
rect 1167 138 1229 150
rect 1167 -138 1183 138
rect 1217 -138 1229 138
rect 1167 -150 1229 -138
<< pdiffc >>
rect -1217 -138 -1183 138
rect -1121 -138 -1087 138
rect -1025 -138 -991 138
rect -929 -138 -895 138
rect -833 -138 -799 138
rect -737 -138 -703 138
rect -641 -138 -607 138
rect -545 -138 -511 138
rect -449 -138 -415 138
rect -353 -138 -319 138
rect -257 -138 -223 138
rect -161 -138 -127 138
rect -65 -138 -31 138
rect 31 -138 65 138
rect 127 -138 161 138
rect 223 -138 257 138
rect 319 -138 353 138
rect 415 -138 449 138
rect 511 -138 545 138
rect 607 -138 641 138
rect 703 -138 737 138
rect 799 -138 833 138
rect 895 -138 929 138
rect 991 -138 1025 138
rect 1087 -138 1121 138
rect 1183 -138 1217 138
<< nsubdiff >>
rect -1297 299 -1235 333
rect 1235 299 1331 333
rect 1297 237 1331 299
rect 1297 -299 1331 -237
<< nsubdiffcont >>
rect -1235 299 1235 333
rect 1297 -237 1331 237
<< poly >>
rect -1167 150 -1137 176
rect -1071 150 -1041 176
rect -975 150 -945 176
rect -879 150 -849 176
rect -783 150 -753 176
rect -687 150 -657 176
rect -591 150 -561 176
rect -495 150 -465 176
rect -399 150 -369 176
rect -303 150 -273 176
rect -207 150 -177 176
rect -111 150 -81 176
rect -15 150 15 176
rect 81 150 111 176
rect 177 150 207 176
rect 273 150 303 176
rect 369 150 399 176
rect 465 150 495 176
rect 561 150 591 176
rect 657 150 687 176
rect 753 150 783 176
rect 849 150 879 176
rect 945 150 975 176
rect 1041 150 1071 176
rect 1137 150 1167 176
rect -1167 -181 -1137 -150
rect -1071 -181 -1041 -150
rect -975 -181 -945 -150
rect -879 -181 -849 -150
rect -783 -181 -753 -150
rect -687 -181 -657 -150
rect -591 -181 -561 -150
rect -495 -181 -465 -150
rect -399 -181 -369 -150
rect -303 -181 -273 -150
rect -207 -181 -177 -150
rect -111 -181 -81 -150
rect -15 -181 15 -150
rect 81 -181 111 -150
rect 177 -181 207 -150
rect 273 -181 303 -150
rect 369 -181 399 -150
rect 465 -181 495 -150
rect 561 -181 591 -150
rect 657 -181 687 -150
rect 753 -181 783 -150
rect 849 -181 879 -150
rect 945 -181 975 -150
rect 1041 -181 1071 -150
rect 1137 -181 1167 -150
rect -1167 -247 1167 -181
<< locali >>
rect -1297 299 -1235 333
rect 1235 299 1331 333
rect 1297 237 1331 299
rect -1217 138 -1183 154
rect -1217 -154 -1183 -138
rect -1121 138 -1087 154
rect -1121 -154 -1087 -138
rect -1025 138 -991 154
rect -1025 -154 -991 -138
rect -929 138 -895 154
rect -929 -154 -895 -138
rect -833 138 -799 154
rect -833 -154 -799 -138
rect -737 138 -703 154
rect -737 -154 -703 -138
rect -641 138 -607 154
rect -641 -154 -607 -138
rect -545 138 -511 154
rect -545 -154 -511 -138
rect -449 138 -415 154
rect -449 -154 -415 -138
rect -353 138 -319 154
rect -353 -154 -319 -138
rect -257 138 -223 154
rect -257 -154 -223 -138
rect -161 138 -127 154
rect -161 -154 -127 -138
rect -65 138 -31 154
rect -65 -154 -31 -138
rect 31 138 65 154
rect 31 -154 65 -138
rect 127 138 161 154
rect 127 -154 161 -138
rect 223 138 257 154
rect 223 -154 257 -138
rect 319 138 353 154
rect 319 -154 353 -138
rect 415 138 449 154
rect 415 -154 449 -138
rect 511 138 545 154
rect 511 -154 545 -138
rect 607 138 641 154
rect 607 -154 641 -138
rect 703 138 737 154
rect 703 -154 737 -138
rect 799 138 833 154
rect 799 -154 833 -138
rect 895 138 929 154
rect 895 -154 929 -138
rect 991 138 1025 154
rect 991 -154 1025 -138
rect 1087 138 1121 154
rect 1087 -154 1121 -138
rect 1183 138 1217 154
rect 1183 -154 1217 -138
rect 1297 -299 1331 -237
<< viali >>
rect -1217 -138 -1183 138
rect -1121 -138 -1087 138
rect -1025 -138 -991 138
rect -929 -138 -895 138
rect -833 -138 -799 138
rect -737 -138 -703 138
rect -641 -138 -607 138
rect -545 -138 -511 138
rect -449 -138 -415 138
rect -353 -138 -319 138
rect -257 -138 -223 138
rect -161 -138 -127 138
rect -65 -138 -31 138
rect 31 -138 65 138
rect 127 -138 161 138
rect 223 -138 257 138
rect 319 -138 353 138
rect 415 -138 449 138
rect 511 -138 545 138
rect 607 -138 641 138
rect 703 -138 737 138
rect 799 -138 833 138
rect 895 -138 929 138
rect 991 -138 1025 138
rect 1087 -138 1121 138
rect 1183 -138 1217 138
<< metal1 >>
rect -1223 138 -1177 150
rect -1223 -138 -1217 138
rect -1183 -138 -1177 138
rect -1223 -150 -1177 -138
rect -1127 138 -1081 150
rect -1127 -138 -1121 138
rect -1087 -138 -1081 138
rect -1127 -150 -1081 -138
rect -1031 138 -985 150
rect -1031 -138 -1025 138
rect -991 -138 -985 138
rect -1031 -150 -985 -138
rect -935 138 -889 150
rect -935 -138 -929 138
rect -895 -138 -889 138
rect -935 -150 -889 -138
rect -839 138 -793 150
rect -839 -138 -833 138
rect -799 -138 -793 138
rect -839 -150 -793 -138
rect -743 138 -697 150
rect -743 -138 -737 138
rect -703 -138 -697 138
rect -743 -150 -697 -138
rect -647 138 -601 150
rect -647 -138 -641 138
rect -607 -138 -601 138
rect -647 -150 -601 -138
rect -551 138 -505 150
rect -551 -138 -545 138
rect -511 -138 -505 138
rect -551 -150 -505 -138
rect -455 138 -409 150
rect -455 -138 -449 138
rect -415 -138 -409 138
rect -455 -150 -409 -138
rect -359 138 -313 150
rect -359 -138 -353 138
rect -319 -138 -313 138
rect -359 -150 -313 -138
rect -263 138 -217 150
rect -263 -138 -257 138
rect -223 -138 -217 138
rect -263 -150 -217 -138
rect -167 138 -121 150
rect -167 -138 -161 138
rect -127 -138 -121 138
rect -167 -150 -121 -138
rect -71 138 -25 150
rect -71 -138 -65 138
rect -31 -138 -25 138
rect -71 -150 -25 -138
rect 25 138 71 150
rect 25 -138 31 138
rect 65 -138 71 138
rect 25 -150 71 -138
rect 121 138 167 150
rect 121 -138 127 138
rect 161 -138 167 138
rect 121 -150 167 -138
rect 217 138 263 150
rect 217 -138 223 138
rect 257 -138 263 138
rect 217 -150 263 -138
rect 313 138 359 150
rect 313 -138 319 138
rect 353 -138 359 138
rect 313 -150 359 -138
rect 409 138 455 150
rect 409 -138 415 138
rect 449 -138 455 138
rect 409 -150 455 -138
rect 505 138 551 150
rect 505 -138 511 138
rect 545 -138 551 138
rect 505 -150 551 -138
rect 601 138 647 150
rect 601 -138 607 138
rect 641 -138 647 138
rect 601 -150 647 -138
rect 697 138 743 150
rect 697 -138 703 138
rect 737 -138 743 138
rect 697 -150 743 -138
rect 793 138 839 150
rect 793 -138 799 138
rect 833 -138 839 138
rect 793 -150 839 -138
rect 889 138 935 150
rect 889 -138 895 138
rect 929 -138 935 138
rect 889 -150 935 -138
rect 985 138 1031 150
rect 985 -138 991 138
rect 1025 -138 1031 138
rect 985 -150 1031 -138
rect 1081 138 1127 150
rect 1081 -138 1087 138
rect 1121 -138 1127 138
rect 1081 -150 1127 -138
rect 1177 138 1223 150
rect 1177 -138 1183 138
rect 1217 -138 1223 138
rect 1177 -150 1223 -138
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1314 -316 1314 316
string parameters w 1.5 l 0.15 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
