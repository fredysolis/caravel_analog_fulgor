magic
tech sky130A
magscale 1 2
timestamp 1624049879
<< isosubstrate >>
rect 17 2892 7722 2988
<< nwell >>
rect 0 2892 7722 2988
rect 2734 996 2771 2154
rect 7685 996 7722 2154
<< pwell >>
rect 1008 774 1054 910
rect 1200 774 1246 910
rect 1392 774 1438 910
rect 1584 774 1630 910
rect 1776 774 1822 910
rect 1968 774 2014 910
rect 2160 774 2206 910
rect 2352 774 2398 910
rect 2544 775 2590 910
rect 6648 570 7722 996
rect 78 0 239 57
rect 0 -96 7722 0
<< psubdiff >>
rect 2630 926 2823 960
rect 6544 926 7686 960
rect 7652 454 7686 926
rect 2630 36 2807 70
rect 4884 36 5058 70
rect 36 -60 132 -26
rect 7590 -60 7614 -26
<< nsubdiff >>
rect 108 2918 132 2952
rect 2602 2918 2866 2952
rect 7590 2918 7614 2952
rect 2630 2822 2808 2856
rect 4884 2822 5058 2856
rect 7652 1066 7686 2258
rect 2804 1032 2887 1066
rect 7581 1032 7686 1066
<< psubdiffcont >>
rect 132 -60 7590 -26
<< nsubdiffcont >>
rect 132 2918 2602 2952
rect 2866 2918 7590 2952
<< poly >>
rect 4929 2641 5056 2661
rect 200 2253 228 2276
rect 2490 2253 2534 2276
rect 200 2210 2534 2253
rect 3216 2084 3540 2342
rect 3894 2276 4788 2347
rect 4929 2300 4950 2641
rect 5034 2342 5056 2641
rect 5034 2300 5363 2342
rect 4929 2276 5363 2300
rect 200 534 2534 544
rect 200 462 220 534
rect 2514 462 2534 534
rect 200 452 2534 462
rect 3222 382 3540 652
rect 4935 452 5061 453
rect 3894 382 4788 448
rect 4935 435 5317 452
rect 4935 243 4957 435
rect 5038 386 5317 435
rect 5038 243 5061 386
rect 4935 222 5061 243
<< polycont >>
rect 228 2253 2490 2299
rect 4950 2300 5034 2641
rect 220 462 2514 534
rect 4957 243 5038 435
<< locali >>
rect 7652 1066 7686 2286
rect 2804 1032 2892 1066
rect 7581 1032 7686 1066
rect 2628 926 2817 960
rect 6542 926 7686 960
rect 204 452 210 544
rect 2524 452 2530 544
rect 7652 450 7686 926
<< viali >>
rect 36 2918 132 2952
rect 132 2918 2602 2952
rect 2602 2918 2866 2952
rect 2866 2918 7590 2952
rect 7590 2918 7686 2952
rect 36 2822 7686 2856
rect 4929 2641 5056 2661
rect 212 2299 2506 2309
rect 212 2253 228 2299
rect 228 2253 2490 2299
rect 2490 2253 2506 2299
rect 4929 2300 4950 2641
rect 4950 2300 5034 2641
rect 5034 2300 5056 2641
rect 4929 2276 5056 2300
rect 212 2243 2506 2253
rect 36 70 70 960
rect 210 534 2524 544
rect 210 462 220 534
rect 220 462 2514 534
rect 2514 462 2524 534
rect 210 452 2524 462
rect 4935 435 5061 453
rect 4935 243 4957 435
rect 4957 243 5038 435
rect 5038 243 5061 435
rect 4935 222 5061 243
rect 36 36 7686 70
rect 36 -60 132 -26
rect 132 -60 7590 -26
rect 7590 -60 7686 -26
<< metal1 >>
rect 0 2952 7722 2958
rect 0 2918 36 2952
rect 7686 2918 7722 2952
rect 0 2856 7722 2918
rect 0 2822 36 2856
rect 7686 2822 7722 2856
rect 0 2816 7722 2822
rect 144 2640 190 2816
rect 336 2616 382 2816
rect 528 2602 574 2816
rect 720 2587 766 2816
rect 912 2596 958 2816
rect 1104 2587 1150 2816
rect 1296 2624 1342 2816
rect 1488 2589 1534 2816
rect 1680 2619 1726 2816
rect 1872 2628 1918 2816
rect 2064 2673 2110 2816
rect 2256 2673 2302 2816
rect 2448 2673 2494 2816
rect 2676 2729 3788 2775
rect 240 2328 286 2420
rect 432 2328 478 2420
rect 624 2328 670 2420
rect 816 2328 862 2420
rect 1008 2328 1054 2420
rect 1200 2328 1246 2420
rect 1392 2328 1438 2420
rect 1584 2328 1630 2420
rect 1776 2328 1822 2420
rect 1968 2328 2014 2420
rect 2160 2328 2206 2420
rect 2352 2328 2398 2420
rect 2544 2328 2590 2518
rect 2676 2328 2780 2729
rect 2974 2673 3020 2729
rect 3166 2673 3212 2729
rect 3358 2673 3404 2729
rect 3550 2673 3596 2729
rect 3742 2673 3788 2729
rect 3934 2673 3980 2816
rect 4126 2673 4172 2816
rect 4318 2673 4364 2816
rect 4510 2673 4556 2816
rect 4702 2673 4748 2816
rect 5132 2673 5178 2816
rect 5324 2673 5370 2816
rect 5516 2673 5562 2816
rect 5708 2673 5754 2816
rect 5900 2673 5946 2816
rect 6092 2673 6138 2816
rect 6284 2673 6330 2816
rect 6476 2673 6522 2816
rect 6668 2673 6714 2816
rect 6860 2673 6906 2816
rect 4923 2661 5062 2673
rect 2865 2385 2875 2661
rect 2927 2385 2937 2661
rect 3057 2385 3067 2661
rect 3119 2385 3129 2661
rect 3249 2385 3259 2661
rect 3311 2385 3321 2661
rect 3441 2385 3451 2661
rect 3503 2385 3513 2661
rect 3633 2385 3643 2661
rect 3695 2385 3705 2661
rect 3825 2385 3835 2661
rect 3887 2385 3897 2661
rect 4017 2385 4027 2661
rect 4079 2385 4089 2661
rect 4209 2385 4219 2661
rect 4271 2385 4281 2661
rect 4401 2385 4411 2661
rect 4463 2385 4473 2661
rect 4593 2385 4603 2661
rect 4655 2385 4665 2661
rect 4785 2385 4795 2661
rect 4847 2385 4856 2661
rect 200 2309 2780 2328
rect 200 2243 212 2309
rect 2506 2243 2780 2309
rect 200 2154 2780 2243
rect 4919 2276 4929 2661
rect 5056 2276 5066 2661
rect 5215 2395 5225 2671
rect 5277 2395 5287 2671
rect 5407 2395 5417 2671
rect 5469 2395 5479 2671
rect 5599 2395 5609 2671
rect 5661 2395 5671 2671
rect 5791 2395 5801 2671
rect 5853 2395 5863 2671
rect 5983 2395 5993 2671
rect 6045 2395 6055 2671
rect 6175 2395 6185 2671
rect 6237 2395 6247 2671
rect 6367 2395 6377 2671
rect 6429 2395 6439 2671
rect 6559 2395 6569 2671
rect 6621 2395 6631 2671
rect 6751 2395 6761 2671
rect 6813 2395 6823 2671
rect 6943 2395 6953 2671
rect 7005 2395 7015 2671
rect 7052 2661 7098 2816
rect 7135 2395 7145 2671
rect 7197 2395 7207 2671
rect 7244 2661 7290 2816
rect 7327 2395 7337 2671
rect 7389 2395 7399 2671
rect 7436 2661 7482 2816
rect 7519 2395 7529 2671
rect 7581 2395 7591 2671
rect 1200 985 1630 2154
rect 4919 1868 5066 2276
rect 2935 1346 7514 1868
rect 0 960 76 972
rect 0 774 36 960
rect 70 774 76 960
rect 240 835 2590 985
rect 240 786 286 835
rect 432 774 478 835
rect 624 774 670 835
rect 817 774 863 835
rect 1008 774 1054 835
rect 1200 774 1246 835
rect 1392 774 1438 835
rect 1584 774 1630 835
rect 1776 774 1822 835
rect 1968 774 2014 835
rect 2160 774 2206 835
rect 2352 774 2398 835
rect 2544 775 2590 835
rect 0 648 10 774
rect 193 648 203 774
rect 322 648 332 774
rect 384 648 394 774
rect 515 648 525 774
rect 577 648 587 774
rect 707 648 717 774
rect 769 648 779 774
rect 899 648 909 774
rect 961 648 971 774
rect 1091 648 1101 774
rect 1153 648 1163 774
rect 1283 648 1293 774
rect 1345 648 1355 774
rect 1475 648 1485 774
rect 1537 648 1547 774
rect 1667 648 1677 774
rect 1729 648 1739 774
rect 1859 648 1869 774
rect 1921 648 1931 774
rect 2051 648 2061 774
rect 2113 648 2123 774
rect 2243 648 2253 774
rect 2305 648 2315 774
rect 2435 648 2445 774
rect 2497 648 2507 774
rect 2878 698 6504 848
rect 0 36 36 648
rect 70 76 76 648
rect 198 544 2780 550
rect 198 452 210 544
rect 2524 452 2780 544
rect 198 446 2780 452
rect 240 360 286 446
rect 432 360 478 446
rect 624 360 670 446
rect 816 360 862 446
rect 1008 360 1054 446
rect 1200 360 1246 446
rect 1392 360 1438 446
rect 1584 360 1630 446
rect 1776 360 1822 446
rect 1968 360 2014 446
rect 2160 360 2206 446
rect 2352 360 2398 446
rect 2544 360 2590 446
rect 144 76 190 223
rect 336 76 382 223
rect 528 76 574 223
rect 720 76 766 224
rect 912 76 958 223
rect 1104 76 1150 223
rect 1296 76 1342 223
rect 1488 76 1534 222
rect 1680 76 1726 223
rect 1872 76 1918 223
rect 2064 76 2110 229
rect 2256 76 2302 230
rect 2448 76 2494 231
rect 2676 165 2780 446
rect 4925 453 5071 698
rect 2865 222 2875 348
rect 2927 222 2937 348
rect 3057 222 3067 348
rect 3119 222 3129 348
rect 3249 222 3259 348
rect 3311 222 3321 348
rect 3441 222 3451 348
rect 3503 222 3513 348
rect 3633 222 3643 348
rect 3695 222 3705 348
rect 3825 222 3835 348
rect 3887 222 3897 348
rect 4017 222 4027 348
rect 4079 222 4089 348
rect 4209 222 4219 348
rect 4271 222 4281 348
rect 4401 222 4411 348
rect 4463 222 4473 348
rect 4593 222 4603 348
rect 4655 222 4665 348
rect 4785 222 4795 348
rect 4847 222 4857 348
rect 4925 222 4935 453
rect 5061 222 5071 453
rect 5215 222 5225 348
rect 5277 222 5287 348
rect 5406 222 5416 348
rect 5468 222 5478 348
rect 5599 222 5609 348
rect 5661 222 5671 348
rect 5791 222 5801 348
rect 5853 222 5863 348
rect 5983 222 5993 348
rect 6045 222 6055 348
rect 6175 222 6185 348
rect 6237 222 6247 348
rect 6367 222 6377 348
rect 6429 222 6439 348
rect 6559 222 6569 348
rect 6621 222 6631 348
rect 6751 222 6761 348
rect 6813 222 6823 348
rect 6943 222 6953 348
rect 7005 222 7015 348
rect 2974 165 3020 212
rect 3166 165 3212 213
rect 3358 165 3404 217
rect 3550 165 3596 217
rect 3742 165 3788 211
rect 2676 119 3788 165
rect 3934 76 3980 211
rect 4126 76 4172 211
rect 4318 76 4364 210
rect 4510 76 4556 211
rect 4702 76 4748 211
rect 4929 210 5067 222
rect 5132 76 5178 217
rect 5324 76 5370 217
rect 5516 76 5562 217
rect 5708 76 5754 218
rect 5900 76 5946 217
rect 6092 76 6138 217
rect 6284 76 6330 217
rect 6476 76 6522 216
rect 6668 76 6714 217
rect 6860 76 6906 217
rect 7052 76 7098 223
rect 7135 222 7145 348
rect 7197 222 7207 348
rect 7244 76 7290 224
rect 7327 222 7337 348
rect 7389 222 7399 348
rect 7436 76 7482 225
rect 7519 222 7529 348
rect 7581 222 7591 348
rect 70 70 7722 76
rect 7686 36 7722 70
rect 0 -26 7722 36
rect 0 -60 36 -26
rect 7686 -60 7722 -26
rect 0 -66 7722 -60
<< via1 >>
rect 2875 2385 2927 2661
rect 3067 2385 3119 2661
rect 3259 2385 3311 2661
rect 3451 2385 3503 2661
rect 3643 2385 3695 2661
rect 3835 2385 3887 2661
rect 4027 2385 4079 2661
rect 4219 2385 4271 2661
rect 4411 2385 4463 2661
rect 4603 2385 4655 2661
rect 4795 2385 4847 2661
rect 4929 2276 5056 2661
rect 5225 2395 5277 2671
rect 5417 2395 5469 2671
rect 5609 2395 5661 2671
rect 5801 2395 5853 2671
rect 5993 2395 6045 2671
rect 6185 2395 6237 2671
rect 6377 2395 6429 2671
rect 6569 2395 6621 2671
rect 6761 2395 6813 2671
rect 6953 2395 7005 2671
rect 7145 2395 7197 2671
rect 7337 2395 7389 2671
rect 7529 2395 7581 2671
rect 10 648 36 774
rect 36 648 70 774
rect 70 648 193 774
rect 332 648 384 774
rect 525 648 577 774
rect 717 648 769 774
rect 909 648 961 774
rect 1101 648 1153 774
rect 1293 648 1345 774
rect 1485 648 1537 774
rect 1677 648 1729 774
rect 1869 648 1921 774
rect 2061 648 2113 774
rect 2253 648 2305 774
rect 2445 648 2497 774
rect 2875 222 2927 348
rect 3067 222 3119 348
rect 3259 222 3311 348
rect 3451 222 3503 348
rect 3643 222 3695 348
rect 3835 222 3887 348
rect 4027 222 4079 348
rect 4219 222 4271 348
rect 4411 222 4463 348
rect 4603 222 4655 348
rect 4795 222 4847 348
rect 4935 222 5061 453
rect 5225 222 5277 348
rect 5416 222 5468 348
rect 5609 222 5661 348
rect 5801 222 5853 348
rect 5993 222 6045 348
rect 6185 222 6237 348
rect 6377 222 6429 348
rect 6569 222 6621 348
rect 6761 222 6813 348
rect 6953 222 7005 348
rect 7145 222 7197 348
rect 7337 222 7389 348
rect 7529 222 7581 348
<< metal2 >>
rect 5225 2671 7581 2681
rect 2875 2661 5056 2671
rect 2927 2385 3067 2661
rect 3119 2385 3259 2661
rect 3311 2385 3451 2661
rect 3503 2385 3643 2661
rect 3695 2385 3835 2661
rect 3887 2385 4027 2661
rect 4079 2385 4219 2661
rect 4271 2385 4411 2661
rect 4463 2385 4603 2661
rect 4655 2385 4795 2661
rect 4847 2385 4929 2661
rect 2875 2375 4929 2385
rect 5277 2395 5417 2671
rect 5469 2395 5609 2671
rect 5661 2395 5801 2671
rect 5853 2395 5993 2671
rect 6045 2395 6185 2671
rect 6237 2395 6377 2671
rect 6429 2395 6569 2671
rect 6621 2395 6761 2671
rect 6813 2395 6953 2671
rect 7005 2395 7145 2671
rect 7197 2395 7337 2671
rect 7389 2395 7529 2671
rect 5225 2385 7581 2395
rect 4929 2266 5056 2276
rect 10 774 2507 784
rect 193 648 332 774
rect 384 648 525 774
rect 577 648 717 774
rect 769 648 909 774
rect 961 648 1101 774
rect 1153 648 1293 774
rect 1345 648 1485 774
rect 1537 648 1677 774
rect 1729 648 1869 774
rect 1921 648 2061 774
rect 2113 648 2253 774
rect 2305 648 2445 774
rect 2497 648 2507 774
rect 10 638 2507 648
rect 4935 453 5061 463
rect 2875 348 4935 358
rect 2927 222 3067 348
rect 3119 222 3259 348
rect 3311 222 3451 348
rect 3503 222 3643 348
rect 3695 222 3835 348
rect 3887 222 4027 348
rect 4079 222 4219 348
rect 4271 222 4411 348
rect 4463 222 4603 348
rect 4655 222 4795 348
rect 4847 222 4935 348
rect 6953 358 7581 2385
rect 2875 212 5061 222
rect 5225 348 7581 358
rect 5277 222 5416 348
rect 5468 222 5609 348
rect 5661 222 5801 348
rect 5853 222 5993 348
rect 6045 222 6185 348
rect 6237 222 6377 348
rect 6429 222 6569 348
rect 6621 222 6761 348
rect 6813 222 6953 348
rect 7005 222 7145 348
rect 7197 222 7337 348
rect 7389 222 7529 348
rect 5225 212 7581 222
use sky130_fd_pr__nfet_01v8_8GRULZ  sky130_fd_pr__nfet_01v8_8GRULZ_0
timestamp 1624049879
transform 1 0 4691 0 1 742
box -1957 -254 1957 254
use sky130_fd_pr__nfet_01v8_MUHGM9  sky130_fd_pr__nfet_01v8_MUHGM9_0
timestamp 1624049879
transform 1 0 3861 0 1 285
box -1127 -285 1127 285
use sky130_fd_pr__nfet_01v8_YCGG98  sky130_fd_pr__nfet_01v8_YCGG98_0
timestamp 1624049879
transform 1 0 6355 0 1 285
box -1367 -285 1367 285
use sky130_fd_pr__pfet_01v8_4ML9WA  sky130_fd_pr__pfet_01v8_4ML9WA_0
timestamp 1624049879
transform 1 0 5228 0 1 1630
box -2457 -634 2457 634
use sky130_fd_pr__nfet_01v8_YCGG98  sky130_fd_pr__nfet_01v8_YCGG98_1
timestamp 1624049879
transform -1 0 1367 0 1 285
box -1367 -285 1367 285
use sky130_fd_pr__nfet_01v8_YCGG98  sky130_fd_pr__nfet_01v8_YCGG98_2
timestamp 1624049879
transform -1 0 1367 0 -1 711
box -1367 -285 1367 285
use sky130_fd_pr__pfet_01v8_ND88ZC  sky130_fd_pr__pfet_01v8_ND88ZC_1
timestamp 1624049879
transform -1 0 1367 0 1 2523
box -1367 -369 1367 369
use sky130_fd_pr__pfet_01v8_ND88ZC  sky130_fd_pr__pfet_01v8_ND88ZC_0
timestamp 1624049879
transform 1 0 6355 0 1 2523
box -1367 -369 1367 369
use sky130_fd_pr__pfet_01v8_NKZXKB  sky130_fd_pr__pfet_01v8_NKZXKB_0
timestamp 1624049879
transform 1 0 3861 0 1 2523
box -1127 -369 1127 369
<< labels >>
rlabel metal2 4957 243 5038 435 1 nswitch
rlabel metal2 4950 2300 5034 2641 1 pswitch
rlabel poly 3222 382 3540 652 1 Down
rlabel metal2 6953 348 7581 2395 1 out
rlabel poly 3894 382 4788 448 1 nDown
rlabel poly 3894 2276 4788 2347 1 Up
rlabel metal1 2676 2224 2780 2775 1 biasp
rlabel metal1 0 2856 7722 2918 1 vdd
rlabel metal1 0 -26 7722 36 1 vss
rlabel metal1 210 452 2524 544 1 iref
rlabel poly 3216 2084 3540 2342 1 nUp
<< end >>
