magic
tech sky130A
magscale 1 2
timestamp 1623449341
<< nwell >>
rect -263 -264 263 264
<< pmos >>
rect -63 -45 -33 45
rect 33 -45 63 45
<< pdiff >>
rect -125 33 -63 45
rect -125 -33 -113 33
rect -79 -33 -63 33
rect -125 -45 -63 -33
rect -33 33 33 45
rect -33 -33 -17 33
rect 17 -33 33 33
rect -33 -45 33 -33
rect 63 33 125 45
rect 63 -33 79 33
rect 113 -33 125 33
rect 63 -45 125 -33
<< pdiffc >>
rect -113 -33 -79 33
rect -17 -33 17 33
rect 79 -33 113 33
<< nsubdiff >>
rect -193 194 -131 228
rect 131 194 193 228
<< nsubdiffcont >>
rect -131 194 131 228
<< poly >>
rect -63 45 -33 71
rect 33 45 63 71
rect -63 -105 -33 -45
rect 33 -105 63 -45
<< locali >>
rect -193 194 -131 228
rect 131 194 193 228
rect -113 33 -79 49
rect -113 -49 -79 -33
rect -17 33 17 49
rect -17 -49 17 -33
rect 79 33 113 49
rect 79 -49 113 -33
<< viali >>
rect -113 -33 -79 33
rect -17 -33 17 33
rect 79 -33 113 33
<< metal1 >>
rect -119 33 -73 45
rect -119 -33 -113 33
rect -79 -33 -73 33
rect -119 -45 -73 -33
rect -23 33 23 45
rect -23 -33 -17 33
rect 17 -33 23 33
rect -23 -45 23 -33
rect 73 33 119 45
rect 73 -33 79 33
rect 113 -33 119 33
rect 73 -45 119 -33
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -210 -211 210 211
string parameters w 0.45 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
