magic
tech sky130A
magscale 1 2
timestamp 1623969746
<< nwell >>
rect -887 -319 887 319
<< pmos >>
rect -687 -100 -657 100
rect -591 -100 -561 100
rect -495 -100 -465 100
rect -399 -100 -369 100
rect -303 -100 -273 100
rect -207 -100 -177 100
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
rect 177 -100 207 100
rect 273 -100 303 100
rect 369 -100 399 100
rect 465 -100 495 100
rect 561 -100 591 100
rect 657 -100 687 100
<< pdiff >>
rect -749 88 -687 100
rect -749 -88 -737 88
rect -703 -88 -687 88
rect -749 -100 -687 -88
rect -657 88 -591 100
rect -657 -88 -641 88
rect -607 -88 -591 88
rect -657 -100 -591 -88
rect -561 88 -495 100
rect -561 -88 -545 88
rect -511 -88 -495 88
rect -561 -100 -495 -88
rect -465 88 -399 100
rect -465 -88 -449 88
rect -415 -88 -399 88
rect -465 -100 -399 -88
rect -369 88 -303 100
rect -369 -88 -353 88
rect -319 -88 -303 88
rect -369 -100 -303 -88
rect -273 88 -207 100
rect -273 -88 -257 88
rect -223 -88 -207 88
rect -273 -100 -207 -88
rect -177 88 -111 100
rect -177 -88 -161 88
rect -127 -88 -111 88
rect -177 -100 -111 -88
rect -81 88 -15 100
rect -81 -88 -65 88
rect -31 -88 -15 88
rect -81 -100 -15 -88
rect 15 88 81 100
rect 15 -88 31 88
rect 65 -88 81 88
rect 15 -100 81 -88
rect 111 88 177 100
rect 111 -88 127 88
rect 161 -88 177 88
rect 111 -100 177 -88
rect 207 88 273 100
rect 207 -88 223 88
rect 257 -88 273 88
rect 207 -100 273 -88
rect 303 88 369 100
rect 303 -88 319 88
rect 353 -88 369 88
rect 303 -100 369 -88
rect 399 88 465 100
rect 399 -88 415 88
rect 449 -88 465 88
rect 399 -100 465 -88
rect 495 88 561 100
rect 495 -88 511 88
rect 545 -88 561 88
rect 495 -100 561 -88
rect 591 88 657 100
rect 591 -88 607 88
rect 641 -88 657 88
rect 591 -100 657 -88
rect 687 88 749 100
rect 687 -88 703 88
rect 737 -88 749 88
rect 687 -100 749 -88
<< pdiffc >>
rect -737 -88 -703 88
rect -641 -88 -607 88
rect -545 -88 -511 88
rect -449 -88 -415 88
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
rect 415 -88 449 88
rect 511 -88 545 88
rect 607 -88 641 88
rect 703 -88 737 88
<< nsubdiff >>
rect -851 249 -755 283
rect 755 249 851 283
rect -851 187 -817 249
rect 817 187 851 249
rect -851 -249 -817 -187
rect 817 -249 851 -187
rect -851 -283 -755 -249
rect 755 -283 851 -249
<< nsubdiffcont >>
rect -755 249 755 283
rect -851 -187 -817 187
rect 817 -187 851 187
rect -755 -283 755 -249
<< poly >>
rect -687 100 -657 126
rect -591 100 -561 126
rect -495 100 -465 126
rect -399 100 -369 126
rect -303 100 -273 126
rect -207 100 -177 126
rect -111 100 -81 126
rect -15 100 15 126
rect 81 100 111 126
rect 177 100 207 126
rect 273 100 303 126
rect 369 100 399 126
rect 465 100 495 126
rect 561 100 591 126
rect 657 100 687 126
rect -687 -131 -657 -100
rect -591 -131 -561 -100
rect -495 -131 -465 -100
rect -399 -131 -369 -100
rect -303 -131 -273 -100
rect -207 -131 -177 -100
rect -111 -131 -81 -100
rect -15 -131 15 -100
rect 81 -131 111 -100
rect 177 -131 207 -100
rect 273 -131 303 -100
rect 369 -131 399 -100
rect 465 -131 495 -100
rect 561 -131 591 -100
rect 657 -131 687 -100
rect -705 -147 705 -131
rect -705 -181 -689 -147
rect -655 -181 -593 -147
rect -559 -181 -497 -147
rect -463 -181 -401 -147
rect -367 -181 -305 -147
rect -271 -181 -209 -147
rect -175 -181 -113 -147
rect -79 -181 -17 -147
rect 17 -181 79 -147
rect 113 -181 175 -147
rect 209 -181 271 -147
rect 305 -181 367 -147
rect 401 -181 463 -147
rect 497 -181 559 -147
rect 593 -181 655 -147
rect 689 -181 705 -147
rect -705 -197 705 -181
<< polycont >>
rect -689 -181 -655 -147
rect -593 -181 -559 -147
rect -497 -181 -463 -147
rect -401 -181 -367 -147
rect -305 -181 -271 -147
rect -209 -181 -175 -147
rect -113 -181 -79 -147
rect -17 -181 17 -147
rect 79 -181 113 -147
rect 175 -181 209 -147
rect 271 -181 305 -147
rect 367 -181 401 -147
rect 463 -181 497 -147
rect 559 -181 593 -147
rect 655 -181 689 -147
<< locali >>
rect -851 249 -755 283
rect 755 249 851 283
rect -851 187 -817 249
rect 817 187 851 249
rect -737 88 -703 104
rect -737 -104 -703 -88
rect -641 88 -607 104
rect -641 -104 -607 -88
rect -545 88 -511 104
rect -545 -104 -511 -88
rect -449 88 -415 104
rect -449 -104 -415 -88
rect -353 88 -319 104
rect -353 -104 -319 -88
rect -257 88 -223 104
rect -257 -104 -223 -88
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect 223 88 257 104
rect 223 -104 257 -88
rect 319 88 353 104
rect 319 -104 353 -88
rect 415 88 449 104
rect 415 -104 449 -88
rect 511 88 545 104
rect 511 -104 545 -88
rect 607 88 641 104
rect 607 -104 641 -88
rect 703 88 737 104
rect 703 -104 737 -88
rect -705 -181 -689 -147
rect 689 -181 705 -147
rect -851 -249 -817 -187
rect 817 -249 851 -187
rect -851 -283 -755 -249
rect 755 -283 851 -249
<< viali >>
rect -737 -88 -703 88
rect -641 -88 -607 88
rect -545 -88 -511 88
rect -449 -88 -415 88
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
rect 415 -88 449 88
rect 511 -88 545 88
rect 607 -88 641 88
rect 703 -88 737 88
rect -689 -181 -655 -147
rect -655 -181 -593 -147
rect -593 -181 -559 -147
rect -559 -181 -497 -147
rect -497 -181 -463 -147
rect -463 -181 -401 -147
rect -401 -181 -367 -147
rect -367 -181 -305 -147
rect -305 -181 -271 -147
rect -271 -181 -209 -147
rect -209 -181 -175 -147
rect -175 -181 -113 -147
rect -113 -181 -79 -147
rect -79 -181 -17 -147
rect -17 -181 17 -147
rect 17 -181 79 -147
rect 79 -181 113 -147
rect 113 -181 175 -147
rect 175 -181 209 -147
rect 209 -181 271 -147
rect 271 -181 305 -147
rect 305 -181 367 -147
rect 367 -181 401 -147
rect 401 -181 463 -147
rect 463 -181 497 -147
rect 497 -181 559 -147
rect 559 -181 593 -147
rect 593 -181 655 -147
rect 655 -181 689 -147
<< metal1 >>
rect -743 88 -697 100
rect -743 -88 -737 88
rect -703 -88 -697 88
rect -743 -100 -697 -88
rect -647 88 -601 100
rect -647 -88 -641 88
rect -607 -88 -601 88
rect -647 -100 -601 -88
rect -551 88 -505 100
rect -551 -88 -545 88
rect -511 -88 -505 88
rect -551 -100 -505 -88
rect -455 88 -409 100
rect -455 -88 -449 88
rect -415 -88 -409 88
rect -455 -100 -409 -88
rect -359 88 -313 100
rect -359 -88 -353 88
rect -319 -88 -313 88
rect -359 -100 -313 -88
rect -263 88 -217 100
rect -263 -88 -257 88
rect -223 -88 -217 88
rect -263 -100 -217 -88
rect -167 88 -121 100
rect -167 -88 -161 88
rect -127 -88 -121 88
rect -167 -100 -121 -88
rect -71 88 -25 100
rect -71 -88 -65 88
rect -31 -88 -25 88
rect -71 -100 -25 -88
rect 25 88 71 100
rect 25 -88 31 88
rect 65 -88 71 88
rect 25 -100 71 -88
rect 121 88 167 100
rect 121 -88 127 88
rect 161 -88 167 88
rect 121 -100 167 -88
rect 217 88 263 100
rect 217 -88 223 88
rect 257 -88 263 88
rect 217 -100 263 -88
rect 313 88 359 100
rect 313 -88 319 88
rect 353 -88 359 88
rect 313 -100 359 -88
rect 409 88 455 100
rect 409 -88 415 88
rect 449 -88 455 88
rect 409 -100 455 -88
rect 505 88 551 100
rect 505 -88 511 88
rect 545 -88 551 88
rect 505 -100 551 -88
rect 601 88 647 100
rect 601 -88 607 88
rect 641 -88 647 88
rect 601 -100 647 -88
rect 697 88 743 100
rect 697 -88 703 88
rect 737 -88 743 88
rect 697 -100 743 -88
rect -701 -147 701 -141
rect -701 -181 -689 -147
rect 689 -181 701 -147
rect -701 -187 701 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -834 -266 834 266
string parameters w 1 l 0.15 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
