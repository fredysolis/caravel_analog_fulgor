magic
tech sky130A
magscale 1 2
timestamp 1624113565
<< nwell >>
rect 1027 2742 4581 3209
<< metal1 >>
rect 1027 6031 9953 6158
rect 1027 4628 3874 6031
rect 4025 5420 4056 5449
rect 1273 3943 1304 3972
rect 2752 3927 2762 3983
rect 2818 3927 3107 3983
rect 5484 3567 5494 3772
rect 5619 3567 5629 3772
rect 9765 3236 9953 6031
rect 1027 2742 9563 3217
rect 9630 2759 9953 3236
rect 5483 2212 5493 2417
rect 5618 2212 5628 2417
rect 1229 2011 1260 2040
rect 2752 2001 2762 2057
rect 2818 2001 3051 2057
rect 1037 1300 3899 1356
rect 1027 -47 3884 1300
rect 4021 539 4052 568
rect 9765 -47 9953 2759
rect 1027 -174 9953 -47
<< via1 >>
rect 2762 3927 2818 3983
rect 5494 3567 5619 3772
rect 5493 2212 5618 2417
rect 2762 2001 2818 2057
<< metal2 >>
rect 9270 4026 9956 4233
rect 2762 3983 2818 3993
rect 2762 3917 2818 3927
rect 3743 3772 5158 3932
rect 5494 3772 5619 3782
rect 3743 3727 5494 3772
rect 4953 3567 5494 3727
rect 5494 3557 5619 3567
rect 5493 2417 5618 2427
rect 4952 2257 5493 2417
rect 3742 2212 5493 2257
rect 2762 2057 2818 2067
rect 3742 2052 5157 2212
rect 5493 2202 5618 2212
rect 2762 1991 2818 2001
rect 9270 1751 9956 1958
<< via2 >>
rect 2762 3927 2818 3983
rect 2762 2001 2818 2057
<< metal3 >>
rect 863 4524 2828 4600
rect 2752 3983 2828 4524
rect 2752 3927 2762 3983
rect 2818 3927 2828 3983
rect 2752 3922 2828 3927
rect 2752 2057 2828 2062
rect 2752 2001 2762 2057
rect 2818 2001 2828 2057
rect 2752 1460 2828 2001
rect 863 1384 2828 1460
use source_follower_buff_nmos  source_follower_buff_nmos_1 ~/sky130-mpw2-fulgor/source_follower_buff_nmos/mag
timestamp 1624043228
transform 1 0 3483 0 -1 4622
box 336 -1409 7209 1545
use source_follower_buff_pmos  source_follower_buff_pmos_1 ~/sky130-mpw2-fulgor/source_follower_buff_pmos/mag
timestamp 1624113565
transform 1 0 1078 0 -1 4373
box -51 -311 3503 1296
use source_follower_buff_nmos  source_follower_buff_nmos_0
timestamp 1624043228
transform 1 0 3483 0 1 1362
box 336 -1409 7209 1545
use source_follower_buff_pmos  source_follower_buff_pmos_0
timestamp 1624113565
transform 1 0 1078 0 1 1611
box -51 -311 3503 1296
<< labels >>
rlabel metal3 899 4542 930 4571 1 inp
rlabel metal1 1273 3943 1304 3972 1 iref1
rlabel metal1 4025 5420 4056 5449 1 iref2
rlabel metal2 9881 4111 9912 4140 1 outp
rlabel metal1 9677 3060 9708 3089 1 avss1p8
rlabel metal1 9451 3068 9482 3097 1 avdd1p8
rlabel metal2 9849 1828 9880 1857 1 outn
rlabel metal1 4021 539 4052 568 1 iref4
rlabel metal1 1229 2011 1260 2040 1 iref3
rlabel metal3 895 1410 926 1439 1 inn
<< end >>
