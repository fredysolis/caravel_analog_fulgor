magic
tech sky130A
magscale 1 2
timestamp 1624115960
<< nwell >>
rect 1572 6 4828 915
rect 2386 -596 4828 6
rect 1572 -1234 4828 -596
<< pwell >>
rect 3200 -1325 3622 -1321
rect 1572 -2058 4828 -1325
<< pmos >>
rect 2586 -377 2616 -177
rect 2682 -377 2712 -177
rect 2778 -377 2808 -177
rect 2874 -377 2904 -177
rect 2970 -377 3000 -177
rect 3400 -377 3430 -177
rect 3496 -377 3526 -177
rect 3592 -377 3622 -177
rect 3688 -377 3718 -177
rect 3784 -377 3814 -177
rect 4214 -377 4244 -177
rect 4310 -377 4340 -177
rect 4406 -377 4436 -177
rect 4502 -377 4532 -177
rect 4598 -377 4628 -177
rect 1772 -1015 1802 -815
rect 1868 -1015 1898 -815
rect 1964 -1015 1994 -815
rect 2060 -1015 2090 -815
rect 2156 -1015 2186 -815
rect 2586 -1015 2616 -815
rect 2682 -1015 2712 -815
rect 2778 -1015 2808 -815
rect 2874 -1015 2904 -815
rect 2970 -1015 3000 -815
rect 3400 -1015 3430 -815
rect 3496 -1015 3526 -815
rect 3592 -1015 3622 -815
rect 3688 -1015 3718 -815
rect 3784 -1015 3814 -815
rect 4214 -1015 4244 -815
rect 4310 -1015 4340 -815
rect 4406 -1015 4436 -815
rect 4502 -1015 4532 -815
rect 4598 -1015 4628 -815
<< nmoslvt >>
rect 3396 -1631 3426 -1531
<< ndiff >>
rect 3338 -1543 3396 -1531
rect 3338 -1619 3350 -1543
rect 3384 -1619 3396 -1543
rect 3338 -1631 3396 -1619
rect 3426 -1543 3484 -1531
rect 3426 -1619 3438 -1543
rect 3472 -1619 3484 -1543
rect 3426 -1631 3484 -1619
<< pdiff >>
rect 3747 449 3813 461
rect 3747 273 3763 449
rect 3797 273 3813 449
rect 3747 261 3813 273
rect 3939 449 4005 461
rect 3939 273 3955 449
rect 3989 273 4005 449
rect 3939 261 4005 273
rect 2524 -189 2586 -177
rect 2524 -365 2536 -189
rect 2570 -365 2586 -189
rect 2524 -377 2586 -365
rect 2616 -189 2682 -177
rect 2616 -365 2632 -189
rect 2666 -365 2682 -189
rect 2616 -377 2682 -365
rect 2712 -189 2778 -177
rect 2712 -365 2728 -189
rect 2762 -365 2778 -189
rect 2712 -377 2778 -365
rect 2808 -189 2874 -177
rect 2808 -365 2824 -189
rect 2858 -365 2874 -189
rect 2808 -377 2874 -365
rect 2904 -189 2970 -177
rect 2904 -365 2920 -189
rect 2954 -365 2970 -189
rect 2904 -377 2970 -365
rect 3000 -189 3062 -177
rect 3000 -365 3016 -189
rect 3050 -365 3062 -189
rect 3000 -377 3062 -365
rect 3338 -189 3400 -177
rect 3338 -365 3350 -189
rect 3384 -365 3400 -189
rect 3338 -377 3400 -365
rect 3430 -189 3496 -177
rect 3430 -365 3446 -189
rect 3480 -365 3496 -189
rect 3430 -377 3496 -365
rect 3526 -189 3592 -177
rect 3526 -365 3542 -189
rect 3576 -365 3592 -189
rect 3526 -377 3592 -365
rect 3622 -189 3688 -177
rect 3622 -365 3638 -189
rect 3672 -365 3688 -189
rect 3622 -377 3688 -365
rect 3718 -189 3784 -177
rect 3718 -365 3734 -189
rect 3768 -365 3784 -189
rect 3718 -377 3784 -365
rect 3814 -189 3876 -177
rect 3814 -365 3830 -189
rect 3864 -365 3876 -189
rect 3814 -377 3876 -365
rect 4152 -189 4214 -177
rect 4152 -365 4164 -189
rect 4198 -365 4214 -189
rect 4152 -377 4214 -365
rect 4244 -189 4310 -177
rect 4244 -365 4260 -189
rect 4294 -365 4310 -189
rect 4244 -377 4310 -365
rect 4340 -189 4406 -177
rect 4340 -365 4356 -189
rect 4390 -365 4406 -189
rect 4340 -377 4406 -365
rect 4436 -189 4502 -177
rect 4436 -365 4452 -189
rect 4486 -365 4502 -189
rect 4436 -377 4502 -365
rect 4532 -189 4598 -177
rect 4532 -365 4548 -189
rect 4582 -365 4598 -189
rect 4532 -377 4598 -365
rect 4628 -189 4690 -177
rect 4628 -365 4644 -189
rect 4678 -365 4690 -189
rect 4628 -377 4690 -365
rect 1710 -827 1772 -815
rect 1710 -1003 1722 -827
rect 1756 -1003 1772 -827
rect 1710 -1015 1772 -1003
rect 1802 -827 1868 -815
rect 1802 -1003 1818 -827
rect 1852 -1003 1868 -827
rect 1802 -1015 1868 -1003
rect 1898 -827 1964 -815
rect 1898 -1003 1914 -827
rect 1948 -1003 1964 -827
rect 1898 -1015 1964 -1003
rect 1994 -827 2060 -815
rect 1994 -1003 2010 -827
rect 2044 -1003 2060 -827
rect 1994 -1015 2060 -1003
rect 2090 -827 2156 -815
rect 2090 -1003 2106 -827
rect 2140 -1003 2156 -827
rect 2090 -1015 2156 -1003
rect 2186 -827 2248 -815
rect 2186 -1003 2202 -827
rect 2236 -1003 2248 -827
rect 2186 -1015 2248 -1003
rect 2524 -827 2586 -815
rect 2524 -1003 2536 -827
rect 2570 -1003 2586 -827
rect 2524 -1015 2586 -1003
rect 2616 -827 2682 -815
rect 2616 -1003 2632 -827
rect 2666 -1003 2682 -827
rect 2616 -1015 2682 -1003
rect 2712 -827 2778 -815
rect 2712 -1003 2728 -827
rect 2762 -1003 2778 -827
rect 2712 -1015 2778 -1003
rect 2808 -827 2874 -815
rect 2808 -1003 2824 -827
rect 2858 -1003 2874 -827
rect 2808 -1015 2874 -1003
rect 2904 -827 2970 -815
rect 2904 -1003 2920 -827
rect 2954 -1003 2970 -827
rect 2904 -1015 2970 -1003
rect 3000 -827 3062 -815
rect 3000 -1003 3016 -827
rect 3050 -1003 3062 -827
rect 3000 -1015 3062 -1003
rect 3338 -827 3400 -815
rect 3338 -1003 3350 -827
rect 3384 -1003 3400 -827
rect 3338 -1015 3400 -1003
rect 3430 -827 3496 -815
rect 3430 -1003 3446 -827
rect 3480 -1003 3496 -827
rect 3430 -1015 3496 -1003
rect 3526 -827 3592 -815
rect 3526 -1003 3542 -827
rect 3576 -1003 3592 -827
rect 3526 -1015 3592 -1003
rect 3622 -827 3688 -815
rect 3622 -1003 3638 -827
rect 3672 -1003 3688 -827
rect 3622 -1015 3688 -1003
rect 3718 -827 3784 -815
rect 3718 -1003 3734 -827
rect 3768 -1003 3784 -827
rect 3718 -1015 3784 -1003
rect 3814 -827 3876 -815
rect 3814 -1003 3830 -827
rect 3864 -1003 3876 -827
rect 3814 -1015 3876 -1003
rect 4152 -827 4214 -815
rect 4152 -1003 4164 -827
rect 4198 -1003 4214 -827
rect 4152 -1015 4214 -1003
rect 4244 -827 4310 -815
rect 4244 -1003 4260 -827
rect 4294 -1003 4310 -827
rect 4244 -1015 4310 -1003
rect 4340 -827 4406 -815
rect 4340 -1003 4356 -827
rect 4390 -1003 4406 -827
rect 4340 -1015 4406 -1003
rect 4436 -827 4502 -815
rect 4436 -1003 4452 -827
rect 4486 -1003 4502 -827
rect 4436 -1015 4502 -1003
rect 4532 -827 4598 -815
rect 4532 -1003 4548 -827
rect 4582 -1003 4598 -827
rect 4532 -1015 4598 -1003
rect 4628 -827 4690 -815
rect 4628 -1003 4644 -827
rect 4678 -1003 4690 -827
rect 4628 -1015 4690 -1003
<< ndiffc >>
rect 3350 -1619 3384 -1543
rect 3438 -1619 3472 -1543
<< pdiffc >>
rect 3763 273 3797 449
rect 3955 273 3989 449
rect 2536 -365 2570 -189
rect 2632 -365 2666 -189
rect 2728 -365 2762 -189
rect 2824 -365 2858 -189
rect 2920 -365 2954 -189
rect 3016 -365 3050 -189
rect 3350 -365 3384 -189
rect 3446 -365 3480 -189
rect 3542 -365 3576 -189
rect 3638 -365 3672 -189
rect 3734 -365 3768 -189
rect 3830 -365 3864 -189
rect 4164 -365 4198 -189
rect 4260 -365 4294 -189
rect 4356 -365 4390 -189
rect 4452 -365 4486 -189
rect 4548 -365 4582 -189
rect 4644 -365 4678 -189
rect 1722 -1003 1756 -827
rect 1818 -1003 1852 -827
rect 1914 -1003 1948 -827
rect 2010 -1003 2044 -827
rect 2106 -1003 2140 -827
rect 2202 -1003 2236 -827
rect 2536 -1003 2570 -827
rect 2632 -1003 2666 -827
rect 2728 -1003 2762 -827
rect 2824 -1003 2858 -827
rect 2920 -1003 2954 -827
rect 3016 -1003 3050 -827
rect 3350 -1003 3384 -827
rect 3446 -1003 3480 -827
rect 3542 -1003 3576 -827
rect 3638 -1003 3672 -827
rect 3734 -1003 3768 -827
rect 3830 -1003 3864 -827
rect 4164 -1003 4198 -827
rect 4260 -1003 4294 -827
rect 4356 -1003 4390 -827
rect 4452 -1003 4486 -827
rect 4548 -1003 4582 -827
rect 4644 -1003 4678 -827
<< psubdiff >>
rect 3236 -1391 3332 -1357
rect 3490 -1391 3586 -1357
rect 3236 -1453 3270 -1391
rect 3552 -1453 3586 -1391
rect 3236 -1709 3270 -1647
rect 3552 -1709 3586 -1647
rect 2814 -1743 3332 -1709
rect 3490 -1743 3586 -1709
rect 2814 -1798 3586 -1743
rect 1646 -2011 1670 -1798
rect 4777 -2011 4801 -1798
<< nsubdiff >>
rect 1611 691 1635 879
rect 4763 698 4787 879
rect 4199 691 4787 698
rect 2835 636 4787 691
rect 1624 406 2741 424
rect 1624 115 1662 406
rect 2706 115 2741 406
rect 1624 76 2741 115
rect 4197 94 4787 636
rect 2422 -28 2518 6
rect 3068 -28 3164 6
rect 2422 -90 2456 -28
rect 3130 -90 3164 -28
rect 2422 -526 2456 -464
rect 3130 -526 3164 -464
rect 2422 -560 2518 -526
rect 3068 -560 3164 -526
rect 3236 -28 3332 6
rect 3882 -28 3978 6
rect 3236 -90 3270 -28
rect 3944 -90 3978 -28
rect 3236 -526 3270 -464
rect 3944 -526 3978 -464
rect 3236 -560 3332 -526
rect 3882 -560 3978 -526
rect 4050 -28 4146 6
rect 4696 -28 4792 6
rect 4050 -90 4084 -28
rect 4758 -90 4792 -28
rect 4050 -526 4084 -464
rect 4758 -526 4792 -464
rect 4050 -560 4146 -526
rect 4696 -560 4792 -526
rect 1608 -666 1704 -632
rect 2254 -666 2350 -632
rect 1608 -728 1642 -666
rect 2316 -728 2350 -666
rect 1608 -1164 1642 -1102
rect 2316 -1164 2350 -1102
rect 1608 -1198 1704 -1164
rect 2254 -1198 2350 -1164
rect 2422 -666 2518 -632
rect 3068 -666 3164 -632
rect 2422 -728 2456 -666
rect 3130 -728 3164 -666
rect 2422 -1164 2456 -1102
rect 3130 -1164 3164 -1102
rect 2422 -1198 2518 -1164
rect 3068 -1198 3164 -1164
rect 3236 -666 3332 -632
rect 3882 -666 3978 -632
rect 3236 -728 3270 -666
rect 3944 -728 3978 -666
rect 3236 -1164 3270 -1102
rect 3944 -1164 3978 -1102
rect 3236 -1198 3332 -1164
rect 3882 -1198 3978 -1164
rect 4050 -666 4146 -632
rect 4696 -666 4792 -632
rect 4050 -728 4084 -666
rect 4758 -728 4792 -666
rect 4050 -1164 4084 -1102
rect 4758 -1164 4792 -1102
rect 4050 -1198 4146 -1164
rect 4696 -1198 4792 -1164
<< psubdiffcont >>
rect 3332 -1391 3490 -1357
rect 3236 -1647 3270 -1453
rect 3552 -1647 3586 -1453
rect 3332 -1743 3490 -1709
rect 1670 -2011 4777 -1798
<< nsubdiffcont >>
rect 1635 698 4763 879
rect 1635 691 4199 698
rect 1662 115 2706 406
rect 2518 -28 3068 6
rect 2422 -464 2456 -90
rect 3130 -464 3164 -90
rect 2518 -560 3068 -526
rect 3332 -28 3882 6
rect 3236 -464 3270 -90
rect 3944 -464 3978 -90
rect 3332 -560 3882 -526
rect 4146 -28 4696 6
rect 4050 -464 4084 -90
rect 4758 -464 4792 -90
rect 4146 -560 4696 -526
rect 1704 -666 2254 -632
rect 1608 -1102 1642 -728
rect 2316 -1102 2350 -728
rect 1704 -1198 2254 -1164
rect 2518 -666 3068 -632
rect 2422 -1102 2456 -728
rect 3130 -1102 3164 -728
rect 2518 -1198 3068 -1164
rect 3332 -666 3882 -632
rect 3236 -1102 3270 -728
rect 3944 -1102 3978 -728
rect 3332 -1198 3882 -1164
rect 4146 -666 4696 -632
rect 4050 -1102 4084 -728
rect 4758 -1102 4792 -728
rect 4146 -1198 4696 -1164
<< poly >>
rect 2586 -177 2616 -151
rect 2682 -177 2712 -151
rect 2778 -177 2808 -151
rect 2874 -177 2904 -151
rect 2970 -177 3000 -151
rect 2586 -408 2616 -377
rect 2682 -408 2712 -377
rect 2778 -408 2808 -377
rect 2874 -408 2904 -377
rect 2970 -408 3000 -377
rect 2568 -424 3018 -408
rect 2568 -458 2616 -424
rect 2974 -458 3018 -424
rect 2568 -474 3018 -458
rect 3400 -177 3430 -151
rect 3496 -177 3526 -151
rect 3592 -177 3622 -151
rect 3688 -177 3718 -151
rect 3784 -177 3814 -151
rect 3400 -408 3430 -377
rect 3496 -408 3526 -377
rect 3592 -408 3622 -377
rect 3688 -408 3718 -377
rect 3784 -408 3814 -377
rect 3382 -424 3832 -408
rect 3382 -458 3430 -424
rect 3788 -458 3832 -424
rect 3382 -474 3832 -458
rect 4214 -177 4244 -151
rect 4310 -177 4340 -151
rect 4406 -177 4436 -151
rect 4502 -177 4532 -151
rect 4598 -177 4628 -151
rect 4214 -408 4244 -377
rect 4310 -408 4340 -377
rect 4406 -408 4436 -377
rect 4502 -408 4532 -377
rect 4598 -408 4628 -377
rect 4196 -424 4646 -408
rect 4196 -458 4244 -424
rect 4602 -458 4646 -424
rect 4196 -474 4646 -458
rect 1754 -734 2204 -718
rect 1754 -768 1802 -734
rect 2160 -768 2204 -734
rect 1754 -784 2204 -768
rect 1772 -815 1802 -784
rect 1868 -815 1898 -784
rect 1964 -815 1994 -784
rect 2060 -815 2090 -784
rect 2156 -815 2186 -784
rect 1772 -1041 1802 -1015
rect 1868 -1041 1898 -1015
rect 1964 -1041 1994 -1015
rect 2060 -1041 2090 -1015
rect 2156 -1041 2186 -1015
rect 2568 -734 3018 -718
rect 2568 -768 2616 -734
rect 2974 -768 3018 -734
rect 2568 -784 3018 -768
rect 2586 -815 2616 -784
rect 2682 -815 2712 -784
rect 2778 -815 2808 -784
rect 2874 -815 2904 -784
rect 2970 -815 3000 -784
rect 2586 -1041 2616 -1015
rect 2682 -1041 2712 -1015
rect 2778 -1041 2808 -1015
rect 2874 -1041 2904 -1015
rect 2970 -1041 3000 -1015
rect 3382 -734 3832 -718
rect 3382 -768 3430 -734
rect 3788 -768 3832 -734
rect 3382 -784 3832 -768
rect 3400 -815 3430 -784
rect 3496 -815 3526 -784
rect 3592 -815 3622 -784
rect 3688 -815 3718 -784
rect 3784 -815 3814 -784
rect 3400 -1041 3430 -1015
rect 3496 -1041 3526 -1015
rect 3592 -1041 3622 -1015
rect 3688 -1041 3718 -1015
rect 3784 -1041 3814 -1015
rect 4196 -734 4646 -718
rect 4196 -768 4244 -734
rect 4602 -768 4646 -734
rect 4196 -784 4646 -768
rect 4214 -815 4244 -784
rect 4310 -815 4340 -784
rect 4406 -815 4436 -784
rect 4502 -815 4532 -784
rect 4598 -815 4628 -784
rect 4214 -1041 4244 -1015
rect 4310 -1041 4340 -1015
rect 4406 -1041 4436 -1015
rect 4502 -1041 4532 -1015
rect 4598 -1041 4628 -1015
rect 2956 -1447 3022 -1421
rect 3378 -1459 3444 -1421
rect 3378 -1493 3394 -1459
rect 3428 -1493 3444 -1459
rect 3378 -1509 3444 -1493
rect 3396 -1531 3426 -1509
rect 3396 -1657 3426 -1631
<< polycont >>
rect 2616 -458 2974 -424
rect 3430 -458 3788 -424
rect 4244 -458 4602 -424
rect 1802 -768 2160 -734
rect 2616 -768 2974 -734
rect 3430 -768 3788 -734
rect 4244 -768 4602 -734
rect 3394 -1493 3428 -1459
<< locali >>
rect 1619 691 1635 879
rect 4763 691 4781 879
rect 2835 636 4228 691
rect 3763 449 3797 465
rect 1624 406 2733 424
rect 1624 115 1662 406
rect 2706 115 2733 406
rect 3763 257 3797 273
rect 3955 449 3989 465
rect 3955 257 3989 273
rect 4199 145 4228 636
rect 4741 145 4781 691
rect 4199 132 4781 145
rect 4195 116 4781 132
rect 1624 76 2733 115
rect 2422 -28 2518 6
rect 3068 -28 3164 6
rect 2422 -90 2456 -28
rect 3130 -90 3164 -28
rect 2536 -189 2570 -173
rect 2536 -381 2570 -365
rect 2632 -189 2666 -173
rect 2632 -381 2666 -365
rect 2728 -189 2762 -173
rect 2728 -381 2762 -365
rect 2824 -189 2858 -173
rect 2824 -381 2858 -365
rect 2920 -189 2954 -173
rect 2920 -381 2954 -365
rect 3016 -189 3050 -173
rect 3016 -381 3050 -365
rect 2587 -458 2616 -424
rect 2974 -458 2999 -424
rect 2422 -526 2456 -464
rect 3130 -526 3164 -464
rect 2422 -560 2518 -526
rect 3068 -560 3164 -526
rect 3236 -28 3332 6
rect 3882 -28 3978 6
rect 3236 -90 3270 -28
rect 3944 -90 3978 -28
rect 3350 -189 3384 -173
rect 3350 -381 3384 -365
rect 3446 -189 3480 -173
rect 3446 -381 3480 -365
rect 3542 -189 3576 -173
rect 3542 -381 3576 -365
rect 3638 -189 3672 -173
rect 3638 -381 3672 -365
rect 3734 -189 3768 -173
rect 3734 -381 3768 -365
rect 3830 -189 3864 -173
rect 3830 -381 3864 -365
rect 3401 -458 3430 -424
rect 3788 -458 3813 -424
rect 3236 -526 3270 -464
rect 3944 -526 3978 -464
rect 3236 -560 3332 -526
rect 3882 -560 3978 -526
rect 4050 -28 4146 6
rect 4696 -28 4792 6
rect 4050 -90 4084 -28
rect 4758 -90 4792 -28
rect 4164 -189 4198 -173
rect 4164 -381 4198 -365
rect 4260 -189 4294 -173
rect 4260 -381 4294 -365
rect 4356 -189 4390 -173
rect 4356 -381 4390 -365
rect 4452 -189 4486 -173
rect 4452 -381 4486 -365
rect 4548 -189 4582 -173
rect 4548 -381 4582 -365
rect 4644 -189 4678 -173
rect 4644 -381 4678 -365
rect 4215 -458 4244 -424
rect 4602 -458 4627 -424
rect 4050 -526 4084 -464
rect 4758 -526 4792 -464
rect 4050 -560 4146 -526
rect 4696 -560 4792 -526
rect 1608 -666 1704 -632
rect 2254 -666 2350 -632
rect 1608 -728 1642 -666
rect 2316 -728 2350 -666
rect 1773 -768 1802 -734
rect 2160 -768 2185 -734
rect 1722 -827 1756 -811
rect 1722 -1019 1756 -1003
rect 1818 -827 1852 -811
rect 1818 -1019 1852 -1003
rect 1914 -827 1948 -811
rect 1914 -1019 1948 -1003
rect 2010 -827 2044 -811
rect 2010 -1019 2044 -1003
rect 2106 -827 2140 -811
rect 2106 -1019 2140 -1003
rect 2202 -827 2236 -811
rect 2202 -1019 2236 -1003
rect 1608 -1164 1642 -1102
rect 2316 -1164 2350 -1102
rect 1608 -1198 1704 -1164
rect 2254 -1198 2350 -1164
rect 2422 -666 2518 -632
rect 3068 -666 3164 -632
rect 2422 -728 2456 -666
rect 3130 -728 3164 -666
rect 2587 -768 2616 -734
rect 2974 -768 2999 -734
rect 2536 -827 2570 -811
rect 2536 -1019 2570 -1003
rect 2632 -827 2666 -811
rect 2632 -1019 2666 -1003
rect 2728 -827 2762 -811
rect 2728 -1019 2762 -1003
rect 2824 -827 2858 -811
rect 2824 -1019 2858 -1003
rect 2920 -827 2954 -811
rect 2920 -1019 2954 -1003
rect 3016 -827 3050 -811
rect 3016 -1019 3050 -1003
rect 2422 -1164 2456 -1102
rect 3130 -1164 3164 -1102
rect 2422 -1198 2518 -1164
rect 3068 -1198 3164 -1164
rect 3236 -666 3332 -632
rect 3882 -666 3978 -632
rect 3236 -728 3270 -666
rect 3944 -728 3978 -666
rect 3401 -768 3430 -734
rect 3788 -768 3813 -734
rect 3350 -827 3384 -811
rect 3350 -1019 3384 -1003
rect 3446 -827 3480 -811
rect 3446 -1019 3480 -1003
rect 3542 -827 3576 -811
rect 3542 -1019 3576 -1003
rect 3638 -827 3672 -811
rect 3638 -1019 3672 -1003
rect 3734 -827 3768 -811
rect 3734 -1019 3768 -1003
rect 3830 -827 3864 -811
rect 3830 -1019 3864 -1003
rect 3236 -1164 3270 -1102
rect 3944 -1164 3978 -1102
rect 3236 -1198 3332 -1164
rect 3882 -1198 3978 -1164
rect 4050 -666 4146 -632
rect 4696 -666 4792 -632
rect 4050 -728 4084 -666
rect 4758 -728 4792 -666
rect 4215 -768 4244 -734
rect 4602 -768 4627 -734
rect 4164 -827 4198 -811
rect 4164 -1019 4198 -1003
rect 4260 -827 4294 -811
rect 4260 -1019 4294 -1003
rect 4356 -827 4390 -811
rect 4356 -1019 4390 -1003
rect 4452 -827 4486 -811
rect 4452 -1019 4486 -1003
rect 4548 -827 4582 -811
rect 4548 -1019 4582 -1003
rect 4644 -827 4678 -811
rect 4644 -1019 4678 -1003
rect 4050 -1164 4084 -1102
rect 4758 -1164 4792 -1102
rect 4050 -1198 4146 -1164
rect 4696 -1198 4792 -1164
rect 3236 -1391 3332 -1357
rect 3490 -1391 3586 -1357
rect 3236 -1453 3270 -1391
rect 3552 -1453 3586 -1391
rect 3378 -1493 3394 -1459
rect 3428 -1493 3444 -1459
rect 3350 -1543 3384 -1527
rect 3350 -1635 3384 -1619
rect 3438 -1543 3472 -1527
rect 3438 -1635 3472 -1619
rect 3236 -1709 3270 -1647
rect 3552 -1709 3586 -1647
rect 2814 -1743 3332 -1709
rect 3490 -1743 3586 -1709
rect 2814 -1798 3586 -1743
rect 1654 -2011 1670 -1798
rect 4777 -2011 4793 -1798
<< viali >>
rect 2592 698 4763 879
rect 2592 691 4199 698
rect 4199 691 4763 698
rect 1662 115 2706 406
rect 3763 273 3797 449
rect 3955 273 3989 449
rect 4228 145 4741 691
rect 2536 -365 2570 -189
rect 2632 -365 2666 -189
rect 2728 -365 2762 -189
rect 2824 -365 2858 -189
rect 2920 -365 2954 -189
rect 3016 -365 3050 -189
rect 2616 -458 2974 -424
rect 3350 -365 3384 -189
rect 3446 -365 3480 -189
rect 3542 -365 3576 -189
rect 3638 -365 3672 -189
rect 3734 -365 3768 -189
rect 3830 -365 3864 -189
rect 3430 -458 3788 -424
rect 4164 -365 4198 -189
rect 4260 -365 4294 -189
rect 4356 -365 4390 -189
rect 4452 -365 4486 -189
rect 4548 -365 4582 -189
rect 4644 -365 4678 -189
rect 4244 -458 4602 -424
rect 1802 -768 2160 -734
rect 1722 -1003 1756 -827
rect 1818 -1003 1852 -827
rect 1914 -1003 1948 -827
rect 2010 -1003 2044 -827
rect 2106 -1003 2140 -827
rect 2202 -1003 2236 -827
rect 2616 -768 2974 -734
rect 2536 -1003 2570 -827
rect 2632 -1003 2666 -827
rect 2728 -1003 2762 -827
rect 2824 -1003 2858 -827
rect 2920 -1003 2954 -827
rect 3016 -1003 3050 -827
rect 3430 -768 3788 -734
rect 3350 -1003 3384 -827
rect 3446 -1003 3480 -827
rect 3542 -1003 3576 -827
rect 3638 -1003 3672 -827
rect 3734 -1003 3768 -827
rect 3830 -1003 3864 -827
rect 4244 -768 4602 -734
rect 4164 -1003 4198 -827
rect 4260 -1003 4294 -827
rect 4356 -1003 4390 -827
rect 4452 -1003 4486 -827
rect 4548 -1003 4582 -827
rect 4644 -1003 4678 -827
rect 2972 -1493 3006 -1425
rect 3394 -1459 3428 -1425
rect 3394 -1493 3428 -1459
rect 3350 -1619 3384 -1543
rect 3438 -1619 3472 -1543
rect 1670 -2011 4777 -1798
<< metal1 >>
rect 1623 879 4775 885
rect 1623 691 1635 879
rect 4763 691 4775 879
rect 1623 685 4228 691
rect 2996 515 3006 570
rect 3405 515 3415 570
rect 3795 514 3805 589
rect 4054 514 4064 589
rect 1650 406 2718 412
rect 1650 115 1662 406
rect 2706 115 2718 406
rect 1650 109 2718 115
rect 2943 42 2989 290
rect 3026 261 3036 461
rect 3088 261 3098 461
rect 3135 42 3181 290
rect 3218 261 3228 461
rect 3280 261 3290 461
rect 3327 42 3373 290
rect 3410 261 3420 461
rect 3472 261 3482 461
rect 3744 261 3754 461
rect 3806 261 3816 461
rect 3853 216 3899 290
rect 3936 261 3946 461
rect 3998 261 4008 461
rect 4045 216 4091 290
rect 4217 216 4228 685
rect 3853 170 4228 216
rect 4217 145 4228 170
rect 4741 685 4775 691
rect 4741 145 4753 685
rect 4875 627 4885 900
rect 5111 627 5121 900
rect 4885 568 5109 627
rect 4875 503 4885 568
rect 5108 503 5118 568
rect 4217 133 4753 145
rect 1706 36 2156 42
rect 1706 -28 1716 36
rect 2146 -28 2156 36
rect 2520 36 3130 42
rect 2520 -28 2530 36
rect 1716 -206 1762 -34
rect 1799 -377 1809 -177
rect 1861 -377 1871 -177
rect 1908 -206 1954 -34
rect 1991 -377 2001 -177
rect 2053 -377 2063 -177
rect 2100 -206 2146 -34
rect 2960 -17 3130 36
rect 2960 -23 2989 -17
rect 2960 -28 2970 -23
rect 2183 -377 2193 -177
rect 2245 -377 2255 -177
rect 2530 -189 2576 -34
rect 2530 -365 2536 -189
rect 2570 -365 2576 -189
rect 2530 -377 2576 -365
rect 2613 -377 2623 -177
rect 2675 -377 2685 -177
rect 2722 -189 2768 -34
rect 2722 -365 2728 -189
rect 2762 -365 2768 -189
rect 2722 -377 2768 -365
rect 2805 -377 2815 -177
rect 2867 -377 2877 -177
rect 2914 -189 2960 -34
rect 3120 -48 3130 -17
rect 3270 36 3784 42
rect 3270 -17 3344 36
rect 3270 -48 3280 -17
rect 3327 -28 3344 -17
rect 3120 -54 3280 -48
rect 3774 -28 3784 36
rect 4148 36 4598 42
rect 4148 -28 4158 36
rect 2914 -365 2920 -189
rect 2954 -365 2960 -189
rect 2914 -377 2960 -365
rect 2997 -377 3007 -177
rect 3059 -377 3069 -177
rect 1908 -424 1954 -418
rect 2594 -424 2993 -418
rect 1770 -476 1780 -424
rect 2179 -476 2189 -424
rect 2584 -476 2594 -424
rect 2993 -476 3003 -424
rect 1908 -716 1954 -476
rect 2100 -716 2146 -476
rect 2722 -716 2768 -476
rect 2914 -716 2960 -476
rect 1770 -734 2189 -716
rect 1770 -768 1802 -734
rect 2160 -768 2189 -734
rect 2584 -734 3003 -716
rect 2584 -768 2616 -734
rect 2974 -768 3003 -734
rect 1780 -774 2179 -768
rect 2594 -774 2993 -768
rect 1716 -827 1762 -815
rect 1716 -1003 1722 -827
rect 1756 -1003 1762 -827
rect 1716 -1158 1762 -1003
rect 1799 -1015 1809 -815
rect 1861 -1015 1871 -815
rect 1908 -827 1954 -815
rect 1908 -1003 1914 -827
rect 1948 -1003 1954 -827
rect 1908 -1158 1954 -1003
rect 1991 -1015 2001 -815
rect 2053 -1015 2063 -815
rect 2100 -827 2146 -815
rect 2100 -1003 2106 -827
rect 2140 -1003 2146 -827
rect 2100 -1158 2146 -1003
rect 2183 -1015 2193 -815
rect 2245 -1015 2255 -815
rect 2530 -827 2576 -815
rect 2530 -1003 2536 -827
rect 2570 -1003 2576 -827
rect 1706 -1228 1716 -1164
rect 2530 -1158 2576 -1003
rect 2613 -1015 2623 -815
rect 2675 -1015 2685 -815
rect 2722 -827 2768 -815
rect 2722 -1003 2728 -827
rect 2762 -1003 2768 -827
rect 2722 -1158 2768 -1003
rect 2805 -1015 2815 -815
rect 2867 -1015 2877 -815
rect 2914 -827 2960 -815
rect 2914 -1003 2920 -827
rect 2954 -1003 2960 -827
rect 2914 -1158 2960 -1003
rect 2997 -1015 3007 -815
rect 3059 -1015 3069 -815
rect 3130 -1138 3270 -54
rect 3344 -189 3390 -34
rect 3344 -365 3350 -189
rect 3384 -365 3390 -189
rect 3344 -377 3390 -365
rect 3427 -377 3437 -177
rect 3489 -377 3499 -177
rect 3536 -189 3582 -34
rect 3536 -365 3542 -189
rect 3576 -365 3582 -189
rect 3536 -377 3582 -365
rect 3619 -377 3629 -177
rect 3681 -377 3691 -177
rect 3728 -189 3774 -34
rect 4588 -28 4598 36
rect 3728 -365 3734 -189
rect 3768 -365 3774 -189
rect 3728 -377 3774 -365
rect 3811 -377 3821 -177
rect 3873 -377 3883 -177
rect 4158 -189 4204 -34
rect 4158 -365 4164 -189
rect 4198 -365 4204 -189
rect 4158 -377 4204 -365
rect 4241 -377 4251 -177
rect 4303 -377 4313 -177
rect 4350 -189 4396 -34
rect 4350 -365 4356 -189
rect 4390 -365 4396 -189
rect 4350 -377 4396 -365
rect 4433 -377 4443 -177
rect 4495 -377 4505 -177
rect 4542 -189 4588 -34
rect 4542 -365 4548 -189
rect 4582 -365 4588 -189
rect 4542 -377 4588 -365
rect 4625 -377 4635 -177
rect 4687 -377 4697 -177
rect 3408 -424 3807 -418
rect 4222 -424 4621 -418
rect 3398 -458 3430 -424
rect 3788 -458 3817 -424
rect 3398 -476 3817 -458
rect 4212 -458 4244 -424
rect 4602 -458 4631 -424
rect 4212 -476 4631 -458
rect 3536 -716 3582 -476
rect 3728 -716 3774 -476
rect 4350 -716 4396 -476
rect 4542 -716 4588 -476
rect 3398 -768 3408 -716
rect 3807 -768 3817 -716
rect 4212 -768 4222 -716
rect 4621 -768 4631 -716
rect 3408 -774 3807 -768
rect 4222 -774 4621 -768
rect 3344 -827 3390 -815
rect 3344 -1003 3350 -827
rect 3384 -1003 3390 -827
rect 2146 -1228 2156 -1164
rect 1706 -1234 2156 -1228
rect 2520 -1228 2530 -1164
rect 3120 -1144 3280 -1138
rect 2960 -1228 2970 -1164
rect 2520 -1234 2970 -1228
rect 3120 -1234 3130 -1144
rect 3270 -1234 3280 -1144
rect 3344 -1158 3390 -1003
rect 3427 -1015 3437 -815
rect 3489 -1015 3499 -815
rect 3536 -827 3582 -815
rect 3536 -1003 3542 -827
rect 3576 -1003 3582 -827
rect 3536 -1158 3582 -1003
rect 3619 -1015 3629 -815
rect 3681 -1015 3691 -815
rect 3728 -827 3774 -815
rect 3728 -1003 3734 -827
rect 3768 -1003 3774 -827
rect 3728 -1158 3774 -1003
rect 3811 -1015 3821 -815
rect 3873 -1015 3883 -815
rect 4158 -827 4204 -815
rect 4158 -1003 4164 -827
rect 4198 -1003 4204 -827
rect 3334 -1228 3344 -1164
rect 4158 -1158 4204 -1003
rect 4241 -1015 4251 -815
rect 4303 -1015 4313 -815
rect 4350 -827 4396 -815
rect 4350 -1003 4356 -827
rect 4390 -1003 4396 -827
rect 4350 -1158 4396 -1003
rect 4433 -1015 4443 -815
rect 4495 -1015 4505 -815
rect 4542 -827 4588 -815
rect 4542 -1003 4548 -827
rect 4582 -1003 4588 -827
rect 4542 -1158 4588 -1003
rect 4625 -1015 4635 -815
rect 4687 -1015 4697 -815
rect 3774 -1228 3784 -1164
rect 3334 -1234 3784 -1228
rect 4148 -1228 4158 -1164
rect 4588 -1228 4598 -1164
rect 4148 -1234 4598 -1228
rect 4885 -1407 5109 503
rect 2952 -1493 2962 -1417
rect 3016 -1493 3026 -1417
rect 3374 -1493 3384 -1417
rect 3438 -1493 3448 -1417
rect 4875 -1459 4885 -1407
rect 5109 -1459 5119 -1407
rect 3382 -1499 3440 -1493
rect 2900 -1631 2910 -1531
rect 3344 -1543 3390 -1531
rect 3010 -1792 3056 -1602
rect 3344 -1619 3350 -1543
rect 3384 -1619 3390 -1543
rect 3344 -1792 3390 -1619
rect 3432 -1631 3438 -1531
rect 3490 -1631 3500 -1531
rect 1658 -1798 4789 -1792
rect 1658 -2011 1670 -1798
rect 4777 -2011 4789 -1798
rect 1658 -2017 4789 -2011
<< via1 >>
rect 1635 691 2592 879
rect 2592 691 4763 879
rect 3006 515 3405 570
rect 3805 514 4054 589
rect 1662 115 2706 406
rect 3036 261 3088 461
rect 3228 261 3280 461
rect 3420 261 3472 461
rect 3754 449 3806 461
rect 3754 273 3763 449
rect 3763 273 3797 449
rect 3797 273 3806 449
rect 3754 261 3806 273
rect 3946 449 3998 461
rect 3946 273 3955 449
rect 3955 273 3989 449
rect 3989 273 3998 449
rect 3946 261 3998 273
rect 4885 627 5111 900
rect 4885 503 5108 568
rect 1716 -34 2146 36
rect 1809 -377 1861 -177
rect 2001 -377 2053 -177
rect 2530 -34 2960 36
rect 2193 -377 2245 -177
rect 2623 -189 2675 -177
rect 2623 -365 2632 -189
rect 2632 -365 2666 -189
rect 2666 -365 2675 -189
rect 2623 -377 2675 -365
rect 2815 -189 2867 -177
rect 2815 -365 2824 -189
rect 2824 -365 2858 -189
rect 2858 -365 2867 -189
rect 2815 -377 2867 -365
rect 3130 -48 3270 42
rect 3344 -34 3774 36
rect 3007 -189 3059 -177
rect 3007 -365 3016 -189
rect 3016 -365 3050 -189
rect 3050 -365 3059 -189
rect 3007 -377 3059 -365
rect 1780 -476 2179 -424
rect 2594 -458 2616 -424
rect 2616 -458 2974 -424
rect 2974 -458 2993 -424
rect 2594 -476 2993 -458
rect 1809 -827 1861 -815
rect 1809 -1003 1818 -827
rect 1818 -1003 1852 -827
rect 1852 -1003 1861 -827
rect 1809 -1015 1861 -1003
rect 2001 -827 2053 -815
rect 2001 -1003 2010 -827
rect 2010 -1003 2044 -827
rect 2044 -1003 2053 -827
rect 2001 -1015 2053 -1003
rect 2193 -827 2245 -815
rect 2193 -1003 2202 -827
rect 2202 -1003 2236 -827
rect 2236 -1003 2245 -827
rect 2193 -1015 2245 -1003
rect 1716 -1228 2146 -1158
rect 2623 -827 2675 -815
rect 2623 -1003 2632 -827
rect 2632 -1003 2666 -827
rect 2666 -1003 2675 -827
rect 2623 -1015 2675 -1003
rect 2815 -827 2867 -815
rect 2815 -1003 2824 -827
rect 2824 -1003 2858 -827
rect 2858 -1003 2867 -827
rect 2815 -1015 2867 -1003
rect 3007 -827 3059 -815
rect 3007 -1003 3016 -827
rect 3016 -1003 3050 -827
rect 3050 -1003 3059 -827
rect 3007 -1015 3059 -1003
rect 3437 -189 3489 -177
rect 3437 -365 3446 -189
rect 3446 -365 3480 -189
rect 3480 -365 3489 -189
rect 3437 -377 3489 -365
rect 3629 -189 3681 -177
rect 3629 -365 3638 -189
rect 3638 -365 3672 -189
rect 3672 -365 3681 -189
rect 3629 -377 3681 -365
rect 4158 -34 4588 36
rect 3821 -189 3873 -177
rect 3821 -365 3830 -189
rect 3830 -365 3864 -189
rect 3864 -365 3873 -189
rect 3821 -377 3873 -365
rect 4251 -189 4303 -177
rect 4251 -365 4260 -189
rect 4260 -365 4294 -189
rect 4294 -365 4303 -189
rect 4251 -377 4303 -365
rect 4443 -189 4495 -177
rect 4443 -365 4452 -189
rect 4452 -365 4486 -189
rect 4486 -365 4495 -189
rect 4443 -377 4495 -365
rect 4635 -189 4687 -177
rect 4635 -365 4644 -189
rect 4644 -365 4678 -189
rect 4678 -365 4687 -189
rect 4635 -377 4687 -365
rect 3408 -734 3807 -716
rect 3408 -768 3430 -734
rect 3430 -768 3788 -734
rect 3788 -768 3807 -734
rect 4222 -734 4621 -716
rect 4222 -768 4244 -734
rect 4244 -768 4602 -734
rect 4602 -768 4621 -734
rect 2530 -1228 2960 -1158
rect 3130 -1234 3270 -1144
rect 3437 -827 3489 -815
rect 3437 -1003 3446 -827
rect 3446 -1003 3480 -827
rect 3480 -1003 3489 -827
rect 3437 -1015 3489 -1003
rect 3629 -827 3681 -815
rect 3629 -1003 3638 -827
rect 3638 -1003 3672 -827
rect 3672 -1003 3681 -827
rect 3629 -1015 3681 -1003
rect 3821 -827 3873 -815
rect 3821 -1003 3830 -827
rect 3830 -1003 3864 -827
rect 3864 -1003 3873 -827
rect 3821 -1015 3873 -1003
rect 3344 -1228 3774 -1158
rect 4251 -827 4303 -815
rect 4251 -1003 4260 -827
rect 4260 -1003 4294 -827
rect 4294 -1003 4303 -827
rect 4251 -1015 4303 -1003
rect 4443 -827 4495 -815
rect 4443 -1003 4452 -827
rect 4452 -1003 4486 -827
rect 4486 -1003 4495 -827
rect 4443 -1015 4495 -1003
rect 4635 -827 4687 -815
rect 4635 -1003 4644 -827
rect 4644 -1003 4678 -827
rect 4678 -1003 4687 -827
rect 4635 -1015 4687 -1003
rect 4158 -1228 4588 -1158
rect 2962 -1425 3016 -1417
rect 2962 -1493 2972 -1425
rect 2972 -1493 3006 -1425
rect 3006 -1493 3016 -1425
rect 3384 -1425 3438 -1417
rect 3384 -1493 3394 -1425
rect 3394 -1493 3428 -1425
rect 3428 -1493 3438 -1425
rect 4885 -1459 5109 -1407
rect 2910 -1631 2962 -1531
rect 3438 -1543 3490 -1531
rect 3438 -1619 3472 -1543
rect 3472 -1619 3490 -1543
rect 3438 -1631 3490 -1619
rect 1670 -2011 4777 -1798
<< metal2 >>
rect 4885 900 5111 910
rect 1635 879 4763 889
rect 1635 681 4763 691
rect 4885 617 5111 627
rect 3805 589 4054 599
rect 2169 570 3405 580
rect 2169 515 3006 570
rect 2169 505 3405 515
rect 3804 514 3805 568
rect 4885 568 5108 578
rect 4054 514 4885 568
rect 3804 503 4885 514
rect 4885 493 5108 503
rect 3036 461 3088 471
rect 1662 406 2706 416
rect 3228 461 3280 471
rect 3088 273 3228 449
rect 3036 251 3088 261
rect 3420 461 3472 471
rect 3280 273 3420 449
rect 3228 251 3280 261
rect 3754 461 3806 471
rect 3472 290 3754 430
rect 3420 251 3472 261
rect 3946 461 3998 471
rect 3806 273 3946 449
rect 3754 251 3806 261
rect 3946 251 3998 261
rect 1662 105 2706 115
rect 1716 36 3130 42
rect 2146 -34 2530 36
rect 2960 -34 3130 36
rect 1716 -40 3130 -34
rect 3120 -48 3130 -40
rect 3270 36 4588 42
rect 3270 -34 3344 36
rect 3774 -34 4158 36
rect 3270 -40 4588 -34
rect 3270 -48 3280 -40
rect 3120 -54 3280 -48
rect 1807 -177 1863 -167
rect 1807 -387 1863 -377
rect 1999 -177 2055 -167
rect 1999 -387 2055 -377
rect 2191 -177 2247 -167
rect 2191 -387 2247 -377
rect 2621 -177 2677 -167
rect 2621 -387 2677 -377
rect 2813 -177 2869 -167
rect 2813 -387 2869 -377
rect 3005 -177 3061 -167
rect 3005 -387 3061 -377
rect 3435 -177 3491 -167
rect 3435 -387 3491 -377
rect 3627 -177 3683 -167
rect 3627 -387 3683 -377
rect 3819 -177 3875 -167
rect 3819 -387 3875 -377
rect 4249 -177 4305 -167
rect 4249 -387 4305 -377
rect 4441 -177 4497 -167
rect 4441 -387 4497 -377
rect 4633 -177 4689 -167
rect 4633 -387 4689 -377
rect 1054 -424 4624 -418
rect 1054 -476 1780 -424
rect 2179 -476 2594 -424
rect 2993 -476 4624 -424
rect 1054 -486 4624 -476
rect 1054 -716 4624 -706
rect 1054 -768 3408 -716
rect 3807 -768 4222 -716
rect 4621 -768 4624 -716
rect 1054 -774 4624 -768
rect 1807 -815 1863 -805
rect 1807 -1025 1863 -1015
rect 1999 -815 2055 -805
rect 1999 -1025 2055 -1015
rect 2191 -815 2247 -805
rect 2191 -1025 2247 -1015
rect 2621 -815 2677 -805
rect 2621 -1025 2677 -1015
rect 2813 -815 2869 -805
rect 2813 -1025 2869 -1015
rect 3005 -815 3061 -805
rect 3005 -1025 3061 -1015
rect 3435 -815 3491 -805
rect 3435 -1025 3491 -1015
rect 3627 -815 3683 -805
rect 3627 -1025 3683 -1015
rect 3819 -815 3875 -805
rect 3819 -1025 3875 -1015
rect 4249 -815 4305 -805
rect 4249 -1025 4305 -1015
rect 4441 -815 4497 -805
rect 4441 -1025 4497 -1015
rect 4633 -815 4689 -805
rect 4633 -1025 4689 -1015
rect 3120 -1144 3280 -1138
rect 3120 -1152 3130 -1144
rect 1716 -1158 3130 -1152
rect 2146 -1228 2530 -1158
rect 2960 -1228 3130 -1158
rect 1716 -1234 3130 -1228
rect 3270 -1152 3280 -1144
rect 3270 -1158 4588 -1152
rect 3270 -1228 3344 -1158
rect 3774 -1228 4158 -1158
rect 3270 -1234 4588 -1228
rect 4885 -1407 5109 -1397
rect 2396 -1417 4885 -1407
rect 2396 -1459 2962 -1417
rect 3016 -1459 3384 -1417
rect 2962 -1503 3016 -1493
rect 3438 -1459 4885 -1417
rect 4885 -1469 5109 -1459
rect 3384 -1503 3438 -1493
rect 2564 -1521 2640 -1511
rect 3760 -1521 3836 -1511
rect 2640 -1631 2910 -1531
rect 2962 -1631 2968 -1531
rect 2640 -1641 2968 -1631
rect 3432 -1631 3438 -1531
rect 3490 -1631 3760 -1531
rect 3432 -1641 3760 -1631
rect 2564 -1651 2640 -1641
rect 3760 -1651 3836 -1641
rect 1670 -1798 4777 -1788
rect 1670 -2021 4777 -2011
<< via2 >>
rect 2592 691 4763 879
rect 4885 627 5111 900
rect 1662 115 2706 406
rect 1807 -377 1809 -177
rect 1809 -377 1861 -177
rect 1861 -377 1863 -177
rect 1999 -377 2001 -177
rect 2001 -377 2053 -177
rect 2053 -377 2055 -177
rect 2191 -377 2193 -177
rect 2193 -377 2245 -177
rect 2245 -377 2247 -177
rect 2621 -377 2623 -177
rect 2623 -377 2675 -177
rect 2675 -377 2677 -177
rect 2813 -377 2815 -177
rect 2815 -377 2867 -177
rect 2867 -377 2869 -177
rect 3005 -377 3007 -177
rect 3007 -377 3059 -177
rect 3059 -377 3061 -177
rect 3435 -377 3437 -177
rect 3437 -377 3489 -177
rect 3489 -377 3491 -177
rect 3627 -377 3629 -177
rect 3629 -377 3681 -177
rect 3681 -377 3683 -177
rect 3819 -377 3821 -177
rect 3821 -377 3873 -177
rect 3873 -377 3875 -177
rect 4249 -377 4251 -177
rect 4251 -377 4303 -177
rect 4303 -377 4305 -177
rect 4441 -377 4443 -177
rect 4443 -377 4495 -177
rect 4495 -377 4497 -177
rect 4633 -377 4635 -177
rect 4635 -377 4687 -177
rect 4687 -377 4689 -177
rect 1807 -1015 1809 -815
rect 1809 -1015 1861 -815
rect 1861 -1015 1863 -815
rect 1999 -1015 2001 -815
rect 2001 -1015 2053 -815
rect 2053 -1015 2055 -815
rect 2191 -1015 2193 -815
rect 2193 -1015 2245 -815
rect 2245 -1015 2247 -815
rect 2621 -1015 2623 -815
rect 2623 -1015 2675 -815
rect 2675 -1015 2677 -815
rect 2813 -1015 2815 -815
rect 2815 -1015 2867 -815
rect 2867 -1015 2869 -815
rect 3005 -1015 3007 -815
rect 3007 -1015 3059 -815
rect 3059 -1015 3061 -815
rect 3435 -1015 3437 -815
rect 3437 -1015 3489 -815
rect 3489 -1015 3491 -815
rect 3627 -1015 3629 -815
rect 3629 -1015 3681 -815
rect 3681 -1015 3683 -815
rect 3819 -1015 3821 -815
rect 3821 -1015 3873 -815
rect 3873 -1015 3875 -815
rect 4249 -1015 4251 -815
rect 4251 -1015 4303 -815
rect 4303 -1015 4305 -815
rect 4441 -1015 4443 -815
rect 4443 -1015 4495 -815
rect 4495 -1015 4497 -815
rect 4633 -1015 4635 -815
rect 4635 -1015 4687 -815
rect 4687 -1015 4689 -815
rect 2564 -1641 2640 -1521
rect 3760 -1641 3836 -1521
rect 1670 -2011 4777 -1798
<< metal3 >>
rect 4875 900 5121 905
rect 1625 879 4773 884
rect 1625 691 2592 879
rect 4763 691 4773 879
rect 1625 686 4773 691
rect 4875 627 4885 900
rect 5111 627 5121 900
rect 4875 622 5121 627
rect 1652 406 2716 411
rect 1652 115 1662 406
rect 2706 115 2716 406
rect 1652 110 2716 115
rect 1797 -177 1873 -172
rect 1989 -177 2065 -172
rect 2181 -177 2257 -172
rect 2611 -177 2687 -172
rect 2803 -177 2879 -172
rect 2995 -177 3071 -172
rect 3425 -177 3501 -172
rect 1793 -377 1803 -177
rect 1867 -377 1877 -177
rect 1985 -377 1995 -177
rect 2059 -377 2069 -177
rect 2177 -377 2187 -177
rect 2251 -377 2261 -177
rect 2607 -377 2617 -177
rect 2681 -377 2691 -177
rect 2799 -377 2809 -177
rect 2873 -377 2883 -177
rect 2991 -377 3001 -177
rect 3065 -377 3075 -177
rect 3425 -377 3435 -177
rect 3491 -377 3501 -177
rect 1797 -815 1873 -377
rect 1797 -1015 1807 -815
rect 1863 -1015 1873 -815
rect 1797 -1122 1873 -1015
rect 1989 -815 2065 -377
rect 1989 -1015 1999 -815
rect 2055 -1015 2065 -815
rect 1989 -1122 2065 -1015
rect 2181 -815 2257 -377
rect 2181 -1015 2191 -815
rect 2247 -1015 2257 -815
rect 2181 -1122 2257 -1015
rect 2611 -815 2687 -377
rect 2611 -1015 2621 -815
rect 2677 -1015 2687 -815
rect 2611 -1122 2687 -1015
rect 2803 -815 2879 -377
rect 2803 -1015 2813 -815
rect 2869 -1015 2879 -815
rect 2803 -1122 2879 -1015
rect 2995 -815 3071 -377
rect 3425 -815 3501 -377
rect 3617 -177 3693 -172
rect 3617 -377 3627 -177
rect 3683 -377 3693 -177
rect 3617 -815 3693 -377
rect 3809 -177 3885 -172
rect 3809 -377 3819 -177
rect 3875 -377 3885 -177
rect 3809 -815 3885 -377
rect 4239 -177 4315 -172
rect 4239 -377 4249 -177
rect 4305 -377 4315 -177
rect 4239 -815 4315 -377
rect 4431 -177 4507 -172
rect 4431 -377 4441 -177
rect 4497 -377 4507 -177
rect 4431 -815 4507 -377
rect 4623 -177 4699 -172
rect 4623 -377 4633 -177
rect 4689 -377 4699 -177
rect 4623 -815 4699 -377
rect 2995 -1015 3005 -815
rect 3061 -1015 3071 -815
rect 3421 -1015 3431 -815
rect 3495 -1015 3505 -815
rect 3613 -1015 3623 -815
rect 3687 -1015 3697 -815
rect 3805 -1015 3815 -815
rect 3879 -1015 3889 -815
rect 4235 -1015 4245 -815
rect 4309 -1015 4319 -815
rect 4427 -1015 4437 -815
rect 4501 -1015 4511 -815
rect 4619 -1015 4629 -815
rect 4693 -1015 4703 -815
rect 2995 -1122 3071 -1015
rect 1797 -1198 3071 -1122
rect 3425 -1122 3501 -1015
rect 3617 -1122 3693 -1015
rect 3809 -1122 3885 -1015
rect 4239 -1122 4315 -1015
rect 4431 -1122 4507 -1015
rect 4623 -1122 4699 -1015
rect 3425 -1198 4699 -1122
rect 2564 -1516 2640 -1198
rect 3760 -1516 3836 -1198
rect 2554 -1521 2650 -1516
rect 2554 -1641 2564 -1521
rect 2640 -1641 2650 -1521
rect 2554 -1646 2650 -1641
rect 3750 -1521 3846 -1516
rect 3750 -1641 3760 -1521
rect 3836 -1641 3846 -1521
rect 3750 -1646 3846 -1641
rect 1660 -1798 4787 -1793
rect 1660 -2011 1670 -1798
rect 4777 -2011 4787 -1798
rect 1660 -2016 4787 -2011
<< via3 >>
rect 2592 691 4763 879
rect 4885 627 5111 900
rect 1803 -377 1807 -177
rect 1807 -377 1863 -177
rect 1863 -377 1867 -177
rect 1995 -377 1999 -177
rect 1999 -377 2055 -177
rect 2055 -377 2059 -177
rect 2187 -377 2191 -177
rect 2191 -377 2247 -177
rect 2247 -377 2251 -177
rect 2617 -377 2621 -177
rect 2621 -377 2677 -177
rect 2677 -377 2681 -177
rect 2809 -377 2813 -177
rect 2813 -377 2869 -177
rect 2869 -377 2873 -177
rect 3001 -377 3005 -177
rect 3005 -377 3061 -177
rect 3061 -377 3065 -177
rect 3431 -1015 3435 -815
rect 3435 -1015 3491 -815
rect 3491 -1015 3495 -815
rect 3623 -1015 3627 -815
rect 3627 -1015 3683 -815
rect 3683 -1015 3687 -815
rect 3815 -1015 3819 -815
rect 3819 -1015 3875 -815
rect 3875 -1015 3879 -815
rect 4245 -1015 4249 -815
rect 4249 -1015 4305 -815
rect 4305 -1015 4309 -815
rect 4437 -1015 4441 -815
rect 4441 -1015 4497 -815
rect 4497 -1015 4501 -815
rect 4629 -1015 4633 -815
rect 4633 -1015 4689 -815
rect 4689 -1015 4693 -815
rect 1670 -2011 4777 -1798
<< metal4 >>
rect 4884 900 5112 901
rect 2564 879 4764 880
rect 2564 691 2592 879
rect 4763 691 4764 879
rect 2564 690 4764 691
rect 4884 627 4885 900
rect 5111 627 5112 900
rect 4884 626 5112 627
rect 1802 -177 5109 -176
rect 1802 -377 1803 -177
rect 1867 -377 1995 -177
rect 2059 -377 2187 -177
rect 2251 -377 2617 -177
rect 2681 -377 2809 -177
rect 2873 -377 3001 -177
rect 3065 -377 5109 -177
rect 1802 -378 5109 -377
rect 1799 -815 5109 -814
rect 1799 -1015 3431 -815
rect 3495 -1015 3623 -815
rect 3687 -1015 3815 -815
rect 3879 -1015 4245 -815
rect 4309 -1015 4437 -815
rect 4501 -1015 4629 -815
rect 4693 -1015 5109 -815
rect 1799 -1016 5109 -1015
rect 1669 -1798 4778 -1797
rect 1669 -2011 1670 -1798
rect 4777 -2011 4778 -1798
rect 1669 -2012 4778 -2011
use sky130_fd_pr__pfet_01v8_2XUYGK  sky130_fd_pr__pfet_01v8_2XUYGK_5
timestamp 1623947381
transform 1 0 1979 0 1 -915
box -407 -319 407 319
use sky130_fd_pr__pfet_01v8_2XUYGK  sky130_fd_pr__pfet_01v8_2XUYGK_6
timestamp 1623947381
transform 1 0 2793 0 1 -915
box -407 -319 407 319
use sky130_fd_pr__pfet_01v8_2XUYGK  sky130_fd_pr__pfet_01v8_2XUYGK_7
timestamp 1623947381
transform 1 0 3607 0 1 -915
box -407 -319 407 319
use sky130_fd_pr__nfet_01v8_lvt_2AP43D  sky130_fd_pr__nfet_01v8_lvt_2AP43D_1
timestamp 1623961588
transform -1 0 3411 0 1 -1550
box -211 -229 211 229
use sky130_fd_pr__nfet_01v8_lvt_2AP43D  sky130_fd_pr__nfet_01v8_lvt_2AP43D_0
timestamp 1623961588
transform 1 0 2989 0 1 -1550
box -211 -229 211 229
use sky130_fd_pr__pfet_01v8_2XUYGK  sky130_fd_pr__pfet_01v8_2XUYGK_8
timestamp 1623947381
transform 1 0 4421 0 1 -915
box -407 -319 407 319
use sky130_fd_pr__pfet_01v8_2XUYGK  sky130_fd_pr__pfet_01v8_2XUYGK_1
timestamp 1623947381
transform 1 0 1979 0 -1 -277
box -407 -319 407 319
use sky130_fd_pr__pfet_01v8_2XUYGK  sky130_fd_pr__pfet_01v8_2XUYGK_2
timestamp 1623947381
transform 1 0 2793 0 -1 -277
box -407 -319 407 319
use sky130_fd_pr__pfet_01v8_2XUYGK  sky130_fd_pr__pfet_01v8_2XUYGK_3
timestamp 1623947381
transform 1 0 3607 0 -1 -277
box -407 -319 407 319
use sky130_fd_pr__pfet_01v8_2XUYGK  sky130_fd_pr__pfet_01v8_2XUYGK_4
timestamp 1623947381
transform 1 0 4421 0 -1 -277
box -407 -319 407 319
use sky130_fd_pr__pfet_01v8_2XUYGK  sky130_fd_pr__pfet_01v8_2XUYGK_0
timestamp 1623947381
transform -1 0 3206 0 1 361
box -407 -319 407 319
use sky130_fd_pr__pfet_01v8_2XL9AN  sky130_fd_pr__pfet_01v8_2XL9AN_0
timestamp 1623969232
transform -1 0 3924 0 1 361
box -311 -319 311 319
<< labels >>
rlabel metal4 4907 -378 5109 -176 1 outp
rlabel metal4 4907 -1016 5109 -814 1 outn
rlabel nwell 2821 696 3536 855 1 avdd1p8
rlabel pwell 2830 -1989 3545 -1830 1 avss1p8
rlabel metal4 4899 640 5089 877 1 clk
rlabel metal1 3130 -1144 3270 -48 1 vp
rlabel metal2 1054 -486 1180 -418 1 inn
rlabel metal2 1054 -774 1180 -706 1 inp
rlabel metal2 2177 505 2303 580 1 vctrl
<< end >>
