magic
tech sky130A
magscale 1 2
timestamp 1623610677
<< pwell >>
rect -263 -305 263 305
<< nmos >>
rect -63 -95 -33 95
rect 33 -95 63 95
<< ndiff >>
rect -125 83 -63 95
rect -125 -83 -113 83
rect -79 -83 -63 83
rect -125 -95 -63 -83
rect -33 83 33 95
rect -33 -83 -17 83
rect 17 -83 33 83
rect -33 -95 33 -83
rect 63 83 125 95
rect 63 -83 79 83
rect 113 -83 125 83
rect 63 -95 125 -83
<< ndiffc >>
rect -113 -83 -79 83
rect -17 -83 17 83
rect 79 -83 113 83
<< psubdiff >>
rect -227 173 -193 235
rect -227 -235 -193 -173
rect -227 -269 -168 -235
rect 178 -269 227 -235
<< psubdiffcont >>
rect -227 -173 -193 173
rect -168 -269 178 -235
<< poly >>
rect -63 95 -33 121
rect 33 95 63 121
rect -63 -117 -33 -95
rect 33 -117 63 -95
rect -81 -133 81 -117
rect -81 -167 -65 -133
rect 65 -167 81 -133
rect -81 -183 81 -167
<< polycont >>
rect -65 -167 65 -133
<< locali >>
rect -227 173 -193 235
rect -113 83 -79 99
rect -113 -99 -79 -83
rect -17 83 17 99
rect -17 -99 17 -83
rect 79 83 113 99
rect 79 -99 113 -83
rect -81 -167 -65 -133
rect 65 -167 81 -133
rect -227 -235 -193 -173
rect -227 -269 -168 -235
rect 178 -269 227 -235
<< viali >>
rect -113 -83 -79 83
rect -17 -83 17 83
rect 79 -83 113 83
rect -65 -167 65 -133
<< metal1 >>
rect -119 84 -73 95
rect -132 -85 -122 84
rect -70 -85 -60 84
rect -23 83 23 95
rect 73 84 119 95
rect -23 -83 -17 83
rect 17 -83 23 83
rect -119 -95 -73 -85
rect -23 -95 23 -83
rect 60 -85 70 84
rect 122 -85 132 84
rect 73 -95 119 -85
rect -77 -133 77 -127
rect -77 -167 -65 -133
rect 65 -167 77 -133
rect -77 -173 77 -167
<< via1 >>
rect -122 83 -70 84
rect -122 -83 -113 83
rect -113 -83 -79 83
rect -79 -83 -70 83
rect -122 -85 -70 -83
rect 70 83 122 84
rect 70 -83 79 83
rect 79 -83 113 83
rect 113 -83 122 83
rect 70 -85 122 -83
<< metal2 >>
rect -122 84 -70 94
rect 70 84 122 94
rect -70 -85 70 84
rect -122 -95 -70 -85
rect 70 -95 122 -85
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -210 -252 210 252
string parameters w 0.95 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
