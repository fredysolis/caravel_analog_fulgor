* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_4798MH VSUBS a_81_n156# a_111_n125# a_15_n125# a_n173_n125#
+ w_n311_n344# a_n111_n156# a_n15_n156# a_n81_n125#
X0 a_n81_n125# a_n111_n156# a_n173_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n15_n156# a_n81_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_81_n156# a_15_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_BHR94T a_n15_n151# w_n311_n335# a_81_n151# a_111_n125#
+ a_15_n125# a_n173_n125# a_n111_n151# a_n81_n125#
X0 a_111_n125# a_81_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n15_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
.ends

.subckt trans_gate m1_187_n605# m1_45_n513# vss vdd
Xsky130_fd_pr__pfet_01v8_4798MH_0 vss vss m1_187_n605# m1_45_n513# m1_45_n513# vdd
+ vss vss m1_187_n605# sky130_fd_pr__pfet_01v8_4798MH
Xsky130_fd_pr__nfet_01v8_BHR94T_0 vdd vss vdd m1_187_n605# m1_45_n513# m1_45_n513#
+ vdd m1_187_n605# sky130_fd_pr__nfet_01v8_BHR94T
.ends

.subckt sky130_fd_pr__pfet_01v8_7KT7MH VSUBS a_n111_n186# a_111_n125# a_15_n125# a_n173_n125#
+ w_n311_n344# a_n81_n125#
X0 a_n81_n125# a_n111_n186# a_n173_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_15_n125# a_n111_n186# a_n81_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_111_n125# a_n111_n186# a_15_n125# w_n311_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS6QM w_n311_n335# a_111_n125# a_15_n125# a_n173_n125#
+ a_n111_n151# a_n81_n125#
X0 a_111_n125# a_n111_n151# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n111_n151# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n111_n151# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
.ends

.subckt inverter_cp_x1 in vss out vdd
Xsky130_fd_pr__pfet_01v8_7KT7MH_0 vss in out vdd vdd vdd out sky130_fd_pr__pfet_01v8_7KT7MH
Xsky130_fd_pr__nfet_01v8_2BS6QM_0 vss out vss vss in out sky130_fd_pr__nfet_01v8_2BS6QM
.ends

.subckt clock_inverter vss CLK vdd CLK_d nCLK_d
Xtrans_gate_0 nCLK_d inverter_cp_x1_0/out vss vdd trans_gate
Xinverter_cp_x1_0 CLK vss inverter_cp_x1_0/out vdd inverter_cp_x1
Xinverter_cp_x1_2 inverter_cp_x1_2/in vss CLK_d vdd inverter_cp_x1
Xinverter_cp_x1_1 CLK vss inverter_cp_x1_2/in vdd inverter_cp_x1
.ends

.subckt sky130_fd_pr__pfet_01v8_MJG8BZ VSUBS a_n125_n95# a_63_n95# w_n263_n314# a_n33_n95#
+ a_n63_n192#
X0 a_63_n95# a_n63_n192# a_n33_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n33_n95# a_n63_n192# a_n125_n95# w_n263_n314# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_2BS854 w_n311_n335# a_n129_n213# a_111_n125# a_15_n125#
+ a_n173_n125# a_n81_n125#
X0 a_111_n125# a_n129_n213# a_15_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n81_n125# a_n129_n213# a_n173_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_15_n125# a_n129_n213# a_n81_n125# w_n311_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_KU9PSX a_n125_n95# a_n33_n95# a_n81_n183# w_n263_n305#
X0 a_n33_n95# a_n81_n183# a_n125_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
X1 a_n125_n95# a_n81_n183# a_n33_n95# w_n263_n305# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=950000u l=150000u
.ends

.subckt latch_diff nQ Q vss CLK vdd nD D
Xsky130_fd_pr__pfet_01v8_MJG8BZ_0 vss vdd vdd vdd nQ Q sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__pfet_01v8_MJG8BZ_1 vss vdd vdd vdd Q nQ sky130_fd_pr__pfet_01v8_MJG8BZ
Xsky130_fd_pr__nfet_01v8_2BS854_0 vss CLK vss m1_657_280# m1_657_280# vss sky130_fd_pr__nfet_01v8_2BS854
Xsky130_fd_pr__nfet_01v8_KU9PSX_0 m1_657_280# Q nD vss sky130_fd_pr__nfet_01v8_KU9PSX
Xsky130_fd_pr__nfet_01v8_KU9PSX_1 m1_657_280# nQ D vss sky130_fd_pr__nfet_01v8_KU9PSX
.ends

.subckt DFlipFlop vss nQ Q D vdd CLK nCLK
Xclock_inverter_0 vss D vdd latch_diff_0/D latch_diff_0/nD clock_inverter
Xlatch_diff_0 latch_diff_1/nD latch_diff_1/D vss CLK vdd latch_diff_0/nD latch_diff_0/D
+ latch_diff
Xlatch_diff_1 nQ Q vss nCLK vdd latch_diff_1/nD latch_diff_1/D latch_diff
.ends

.subckt sky130_fd_pr__pfet_01v8_ZP3U9B VSUBS a_n221_n84# a_159_n84# w_n359_n303# a_n63_n110#
+ a_n129_n84# a_33_n110# a_n159_n110# a_63_n84# a_129_n110# a_n33_n84#
X0 a_n129_n84# a_n159_n110# a_n221_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_63_n84# a_33_n110# a_n33_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_n33_n84# a_n63_n110# a_n129_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_159_n84# a_129_n110# a_63_n84# w_n359_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_DXA56D w_n359_n252# a_n33_n42# a_129_n68# a_n159_n68#
+ a_n221_n42# a_159_n42# a_n129_n42# a_33_n68# a_n63_n68# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n129_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_159_n42# a_129_n68# a_63_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_n129_n42# a_n159_n68# a_n221_n42# w_n359_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt inverter_min_x4 vdd in vss out
Xsky130_fd_pr__pfet_01v8_ZP3U9B_0 vss out out vdd in vdd in in vdd in out sky130_fd_pr__pfet_01v8_ZP3U9B
Xsky130_fd_pr__nfet_01v8_DXA56D_0 vss out in in out out vss in in vss sky130_fd_pr__nfet_01v8_DXA56D
.ends

.subckt sky130_fd_pr__pfet_01v8_BDRUME VSUBS a_351_n84# a_n513_n84# a_639_n84# a_159_n84#
+ a_n321_n84# a_447_n84# a_n753_n181# a_n609_n84# w_n935_n303# a_n129_n84# a_735_n84#
+ a_255_n84# a_n417_n84# a_63_n84# a_543_n84# a_n705_n84# a_n225_n84# a_n797_n84#
+ a_n33_n84#
X0 a_n705_n84# a_n753_n181# a_n797_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_n513_n84# a_n753_n181# a_n609_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_n417_n84# a_n753_n181# a_n513_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_n321_n84# a_n753_n181# a_n417_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_n225_n84# a_n753_n181# a_n321_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 a_n129_n84# a_n753_n181# a_n225_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 a_n609_n84# a_n753_n181# a_n705_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_63_n84# a_n753_n181# a_n33_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_n33_n84# a_n753_n181# a_n129_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_159_n84# a_n753_n181# a_63_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_255_n84# a_n753_n181# a_159_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 a_351_n84# a_n753_n181# a_255_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 a_543_n84# a_n753_n181# a_447_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 a_447_n84# a_n753_n181# a_351_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 a_639_n84# a_n753_n181# a_543_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_735_n84# a_n753_n181# a_639_n84# w_n935_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_QQE8KM a_543_n42# a_n705_n42# a_n225_n42# a_n797_n42#
+ a_n33_n42# a_351_n42# a_n513_n42# a_639_n42# a_159_n42# w_n935_n252# a_n757_64#
+ a_n321_n42# a_447_n42# a_n609_n42# a_n129_n42# a_735_n42# a_255_n42# a_n417_n42#
+ a_63_n42#
X0 a_63_n42# a_n757_64# a_n33_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n757_64# a_n129_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_351_n42# a_n757_64# a_255_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_159_n42# a_n757_64# a_63_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_255_n42# a_n757_64# a_159_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_447_n42# a_n757_64# a_351_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_543_n42# a_n757_64# a_447_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_735_n42# a_n757_64# a_639_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_639_n42# a_n757_64# a_543_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_n321_n42# a_n757_64# a_n417_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_n705_n42# a_n757_64# a_n797_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_n513_n42# a_n757_64# a_n609_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_n417_n42# a_n757_64# a_n513_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_n225_n42# a_n757_64# a_n321_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_n129_n42# a_n757_64# a_n225_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_n609_n42# a_n757_64# a_n705_n42# w_n935_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt inverter_min_x16 in out vss vdd
Xsky130_fd_pr__pfet_01v8_BDRUME_0 vss out vdd vdd out vdd vdd in out vdd vdd out vdd
+ out vdd out vdd out out out sky130_fd_pr__pfet_01v8_BDRUME
Xsky130_fd_pr__nfet_01v8_QQE8KM_0 out vss out out out out vss vss out vss in vss vss
+ out vss out vss out vss sky130_fd_pr__nfet_01v8_QQE8KM
.ends

.subckt sky130_fd_pr__pfet_01v8_75PKJG VSUBS a_n33_n102# w_n359_n321# a_n177_n199#
+ a_63_n102# a_n129_n102# a_n221_n102# a_25_n199# a_159_n102#
X0 a_159_n102# a_25_n199# a_63_n102# w_n359_n321# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
X1 a_63_n102# a_25_n199# a_n33_n102# w_n359_n321# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
X2 a_n129_n102# a_n177_n199# a_n221_n102# w_n359_n321# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
X3 a_n33_n102# a_n177_n199# a_n129_n102# w_n359_n321# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_XRJ78J a_n33_n102# w_n263_n312# a_63_n102# a_n125_n102#
+ a_n81_124#
X0 a_n33_n102# a_n81_124# a_n125_n102# w_n263_n312# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
X1 a_63_n102# a_n81_124# a_n33_n102# w_n263_n312# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.02e+06u l=150000u
.ends

.subckt nand_logic avss1p8 in1 avdd1p8 in2 out
Xsky130_fd_pr__pfet_01v8_75PKJG_0 avss1p8 avdd1p8 avdd1p8 in1 out out avdd1p8 in2
+ avdd1p8 sky130_fd_pr__pfet_01v8_75PKJG
Xsky130_fd_pr__nfet_01v8_XRJ78J_0 m1_21_n341# avss1p8 avss1p8 avss1p8 in1 sky130_fd_pr__nfet_01v8_XRJ78J
Xsky130_fd_pr__nfet_01v8_XRJ78J_1 out avss1p8 m1_21_n341# m1_21_n341# in2 sky130_fd_pr__nfet_01v8_XRJ78J
.ends

.subckt res_amp_sync_v2 vss avdd1p8 clk_amp clkn clkp rst
XDFlipFlop_0 vss DFlipFlop_0/nQ DFlipFlop_0/Q DFlipFlop_3/D avdd1p8 clkp clkn DFlipFlop
XDFlipFlop_1 vss DFlipFlop_1/nQ DFlipFlop_2/D DFlipFlop_1/D avdd1p8 DFlipFlop_3/D
+ DFlipFlop_0/Q DFlipFlop
XDFlipFlop_2 vss DFlipFlop_2/nQ DFlipFlop_2/Q DFlipFlop_2/D avdd1p8 clkp clkn DFlipFlop
XDFlipFlop_3 vss DFlipFlop_3/nQ DFlipFlop_3/Q DFlipFlop_3/D avdd1p8 clkp clkn DFlipFlop
Xinverter_min_x4_0 avdd1p8 DFlipFlop_0/Q vss DFlipFlop_3/D inverter_min_x4
Xinverter_min_x4_1 avdd1p8 nand_logic_0/out vss DFlipFlop_4/D inverter_min_x4
XDFlipFlop_4 vss DFlipFlop_4/nQ DFlipFlop_4/Q DFlipFlop_4/D avdd1p8 clkp clkn DFlipFlop
Xinverter_min_x4_2 avdd1p8 DFlipFlop_2/D vss DFlipFlop_1/D inverter_min_x4
Xinverter_min_x4_3 avdd1p8 nand_logic_1/out vss rst inverter_min_x4
Xinverter_min_x4_4 avdd1p8 DFlipFlop_4/Q vss inverter_min_x4_4/out inverter_min_x4
Xinverter_min_x16_0 inverter_min_x4_4/out clk_amp vss avdd1p8 inverter_min_x16
Xnand_logic_0 vss DFlipFlop_2/Q avdd1p8 DFlipFlop_3/Q nand_logic_0/out nand_logic
Xnand_logic_1 vss DFlipFlop_4/D avdd1p8 clkp nand_logic_1/out nand_logic
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_4L9VGG VSUBS a_291_n200# w_n487_n419# a_35_n200#
+ a_n291_n238# a_n93_n200# a_163_n200# a_n349_n200# a_n221_n200#
X0 a_291_n200# a_n291_n238# a_163_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X1 a_n221_n200# a_n291_n238# a_n349_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X2 a_35_n200# a_n291_n238# a_n93_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X3 a_163_n200# a_n291_n238# a_35_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X4 a_n93_n200# a_n291_n238# a_n221_n200# w_n487_n419# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
.ends

.subckt sky130_fd_pr__nfet_01v8_L78GGD a_n73_n73# w_n211_n221# a_15_n73# a_n33_33#
X0 a_15_n73# a_n33_33# a_n73_n73# w_n211_n221# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_6RX2PQ VSUBS w_n211_n268# a_15_n48# a_n33_n145# a_n73_n48#
X0 a_15_n48# a_n33_n145# a_n73_n48# w_n211_n268# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt inverter_min vdd out in vss
XXM1 vss vss out in sky130_fd_pr__nfet_01v8_L78GGD
XXM2 vss vdd out in vdd sky130_fd_pr__pfet_01v8_6RX2PQ
.ends

.subckt buffer_no_inv_x05 VSUBS in avdd1p8 out
Xinverter_min_1 avdd1p8 out inverter_min_1/in VSUBS inverter_min
Xinverter_min_0 avdd1p8 inverter_min_1/in in VSUBS inverter_min
.ends

.subckt sky130_fd_pr__pfet_01v8_XA7ZMQ VSUBS a_21_142# a_63_n111# a_n87_142# a_n125_n111#
+ w_n263_n330# a_n33_n111#
X0 a_n33_n111# a_n87_142# a_n125_n111# w_n263_n330# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.11e+06u l=150000u
X1 a_63_n111# a_21_142# a_n33_n111# w_n263_n330# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.11e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_HAN8QX a_15_n142# a_n33_102# a_n73_n142# w_n211_n290#
X0 a_15_n142# a_n33_102# a_n73_n142# w_n211_n290# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.11e+06u l=150000u
.ends

.subckt mux_2to1_logic sel avdd1p8 w_947_n633# avss1p8 out DinA DinB
Xinverter_min_0 avdd1p8 sel_b sel avss1p8 inverter_min
Xsky130_fd_pr__pfet_01v8_XA7ZMQ_0 avss1p8 sel DinA sel DinA avdd1p8 out sky130_fd_pr__pfet_01v8_XA7ZMQ
Xsky130_fd_pr__pfet_01v8_XA7ZMQ_1 avss1p8 sel_b DinB sel_b DinB avdd1p8 out sky130_fd_pr__pfet_01v8_XA7ZMQ
Xsky130_fd_pr__nfet_01v8_HAN8QX_0 out sel_b DinA avss1p8 sky130_fd_pr__nfet_01v8_HAN8QX
Xsky130_fd_pr__nfet_01v8_HAN8QX_1 out sel DinB avss1p8 sky130_fd_pr__nfet_01v8_HAN8QX
.ends

.subckt delay_cell_buff clk clk_out avss1p8 avdd1p8 reg0 reg2 reg1 mux_2to1_logic_5/w_947_n633#
Xbuffer_no_inv_x05_8 avss1p8 mux_2to1_logic_3/DinA avdd1p8 buffer_no_inv_x05_9/in
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_9 avss1p8 buffer_no_inv_x05_9/in avdd1p8 mux_2to1_logic_3/DinB
+ buffer_no_inv_x05
Xmux_2to1_logic_0 reg2 avdd1p8 mux_2to1_logic_0/w_947_n633# avss1p8 mux_2to1_logic_0/out
+ clk mux_2to1_logic_0/DinB mux_2to1_logic
Xmux_2to1_logic_1 reg2 avdd1p8 mux_2to1_logic_1/w_947_n633# avss1p8 mux_2to1_logic_1/out
+ mux_2to1_logic_1/DinA mux_2to1_logic_1/DinB mux_2to1_logic
Xmux_2to1_logic_2 reg1 avdd1p8 mux_2to1_logic_2/w_947_n633# avss1p8 mux_2to1_logic_2/out
+ mux_2to1_logic_0/out mux_2to1_logic_1/out mux_2to1_logic
Xmux_2to1_logic_3 reg2 avdd1p8 mux_2to1_logic_3/w_947_n633# avss1p8 mux_2to1_logic_3/out
+ mux_2to1_logic_3/DinA mux_2to1_logic_3/DinB mux_2to1_logic
Xmux_2to1_logic_4 reg2 avdd1p8 mux_2to1_logic_4/w_947_n633# avss1p8 mux_2to1_logic_4/out
+ mux_2to1_logic_4/DinA mux_2to1_logic_4/DinB mux_2to1_logic
Xmux_2to1_logic_5 reg1 avdd1p8 mux_2to1_logic_5/w_947_n633# avss1p8 mux_2to1_logic_5/out
+ mux_2to1_logic_3/out mux_2to1_logic_4/out mux_2to1_logic
Xmux_2to1_logic_6 reg0 avdd1p8 mux_2to1_logic_6/w_947_n633# avss1p8 nand_logic_0/in1
+ mux_2to1_logic_2/out mux_2to1_logic_5/out mux_2to1_logic
Xbuffer_no_inv_x05_10 avss1p8 mux_2to1_logic_3/DinB avdd1p8 buffer_no_inv_x05_11/in
+ buffer_no_inv_x05
Xnand_logic_0 avss1p8 nand_logic_0/in1 avdd1p8 clk clk_out nand_logic
Xbuffer_no_inv_x05_11 avss1p8 buffer_no_inv_x05_11/in avdd1p8 mux_2to1_logic_4/DinA
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_12 avss1p8 mux_2to1_logic_4/DinA avdd1p8 buffer_no_inv_x05_13/in
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_13 avss1p8 buffer_no_inv_x05_13/in avdd1p8 mux_2to1_logic_4/DinB
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_0 avss1p8 clk avdd1p8 buffer_no_inv_x05_1/in buffer_no_inv_x05
Xbuffer_no_inv_x05_2 avss1p8 mux_2to1_logic_0/DinB avdd1p8 buffer_no_inv_x05_3/in
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_1 avss1p8 buffer_no_inv_x05_1/in avdd1p8 mux_2to1_logic_0/DinB
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_3 avss1p8 buffer_no_inv_x05_3/in avdd1p8 mux_2to1_logic_1/DinA
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_4 avss1p8 mux_2to1_logic_1/DinA avdd1p8 buffer_no_inv_x05_5/in
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_5 avss1p8 buffer_no_inv_x05_5/in avdd1p8 mux_2to1_logic_1/DinB
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_6 avss1p8 mux_2to1_logic_1/DinB avdd1p8 buffer_no_inv_x05_7/in
+ buffer_no_inv_x05
Xbuffer_no_inv_x05_7 avss1p8 buffer_no_inv_x05_7/in avdd1p8 mux_2to1_logic_3/DinA
+ buffer_no_inv_x05
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_72JNYZ a_n81_n100# w_n311_n310# a_n128_122# a_111_n100#
+ a_15_n100# a_n173_n100#
X0 a_15_n100# a_n128_122# a_n81_n100# w_n311_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n81_n100# a_n128_122# a_n173_n100# w_n311_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_111_n100# a_n128_122# a_15_n100# w_n311_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_2XL9AN VSUBS w_n311_n319# a_n81_n100# a_111_n100#
+ a_n129_131# a_15_n100# a_n173_n100#
X0 a_15_n100# a_n129_131# a_n81_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_n100# a_n129_131# a_15_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n81_n100# a_n129_131# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_2XUYGK VSUBS a_n269_n100# a_n81_n100# w_n407_n319#
+ a_111_n100# a_n177_n100# a_15_n100# a_207_n100# a_n225_131#
X0 a_207_n100# a_n225_131# a_111_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_15_n100# a_n225_131# a_n81_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_111_n100# a_n225_131# a_15_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n81_n100# a_n225_131# a_n177_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n177_n100# a_n225_131# a_n269_n100# w_n407_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_2AP43D a_15_n81# a_n33_41# w_n211_n229# a_n73_n81#
X0 a_15_n81# a_n33_41# a_n73_n81# w_n211_n229# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
.ends

.subckt res_amp_lin clk vctrl avdd1p8 avss1p8 inn outn outp inp
Xsky130_fd_pr__pfet_01v8_2XL9AN_0 avss1p8 avdd1p8 a_3747_261# a_3747_261# clk avdd1p8
+ avdd1p8 sky130_fd_pr__pfet_01v8_2XL9AN
Xsky130_fd_pr__pfet_01v8_2XUYGK_0 avss1p8 a_3747_261# a_3747_261# avdd1p8 a_3747_261#
+ vp vp vp vctrl sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_1 avss1p8 vp vp avdd1p8 vp outp outp outp inn sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__nfet_01v8_lvt_2AP43D_0 avss1p8 clk avss1p8 outp sky130_fd_pr__nfet_01v8_lvt_2AP43D
Xsky130_fd_pr__pfet_01v8_2XUYGK_2 avss1p8 vp vp avdd1p8 vp outp outp outp inn sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__nfet_01v8_lvt_2AP43D_1 avss1p8 clk avss1p8 outn sky130_fd_pr__nfet_01v8_lvt_2AP43D
Xsky130_fd_pr__pfet_01v8_2XUYGK_3 avss1p8 vp vp avdd1p8 vp outn outn outn inp sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_4 avss1p8 vp vp avdd1p8 vp outn outn outn inp sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_5 avss1p8 vp vp avdd1p8 vp outp outp outp inn sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_6 avss1p8 vp vp avdd1p8 vp outp outp outp inn sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_7 avss1p8 vp vp avdd1p8 vp outn outn outn inp sky130_fd_pr__pfet_01v8_2XUYGK
Xsky130_fd_pr__pfet_01v8_2XUYGK_8 avss1p8 vp vp avdd1p8 vp outn outn outn inp sky130_fd_pr__pfet_01v8_2XUYGK
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_595QY5 a_n269_n100# a_n81_n100# a_111_n100# a_n177_n100#
+ a_15_n100# w_n407_n310# a_207_n100# a_n225_n188#
X0 a_207_n100# a_n225_n188# a_111_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_15_n100# a_n225_n188# a_n81_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n81_n100# a_n225_n188# a_n177_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_111_n100# a_n225_n188# a_15_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n177_n100# a_n225_n188# a_n269_n100# w_n407_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_9B2JY7 a_n317_n100# a_n33_n100# a_n225_n100# a_n271_122#
+ a_63_n100# a_n129_n100# w_n455_n310# a_255_n100# a_159_n100#
X0 a_63_n100# a_n271_122# a_n33_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n271_122# a_n129_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_159_n100# a_n271_122# a_63_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_255_n100# a_n271_122# a_159_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n225_n100# a_n271_122# a_n317_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n129_n100# a_n271_122# a_n225_n100# w_n455_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_MVT43V a_n33_n100# w_n263_n310# a_63_n100# a_n79_122#
+ a_n125_n100#
X0 a_63_n100# a_n79_122# a_n33_n100# w_n263_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n79_122# a_n125_n100# w_n263_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_NMSMYT a_n33_n100# a_n321_n100# a_n225_n100# w_n551_n310#
+ a_63_n100# a_n368_122# a_n129_n100# a_351_n100# a_255_n100# a_n413_n100# a_159_n100#
X0 a_63_n100# a_n368_122# a_n33_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n368_122# a_n129_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_159_n100# a_n368_122# a_63_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_255_n100# a_n368_122# a_159_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_351_n100# a_n368_122# a_255_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n321_n100# a_n368_122# a_n413_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n225_n100# a_n368_122# a_n321_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n129_n100# a_n368_122# a_n225_n100# w_n551_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_XAYTAL VSUBS w_n311_n319# a_n81_n100# a_n129_n197#
+ a_111_n100# a_15_n100# a_n173_n100#
X0 a_15_n100# a_n129_n197# a_n81_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_n100# a_n129_n197# a_15_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n81_n100# a_n129_n197# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_B2JNY3 a_n33_n100# a_63_n100# a_n221_n100# a_n129_n100#
+ w_n359_n310# a_n176_122# a_159_n100#
X0 a_63_n100# a_n176_122# a_n33_n100# w_n359_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n176_122# a_n129_n100# w_n359_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_159_n100# a_n176_122# a_63_n100# w_n359_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n129_n100# a_n176_122# a_n221_n100# w_n359_n310# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_XACJHL VSUBS a_n81_n197# w_n263_n319# a_n33_n100#
+ a_63_n100# a_n125_n100#
X0 a_63_n100# a_n81_n197# a_n33_n100# w_n263_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n197# a_n125_n100# w_n263_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt iref_ctrl_res_amp vctrl avdd1p8 reg0 reg1 reg2 iref avss1p8
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_0 iref m1_n356_n363# m1_n356_n363# iref iref iref
+ avss1p8 iref m1_n356_n363# sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_1 avss1p8 m1_n356_n363# m1_n356_n363# avdd1p8
+ avss1p8 avss1p8 avss1p8 avss1p8 m1_n356_n363# sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_MVT43V_0 m1_964_n363# avss1p8 vctrl iref vctrl sky130_fd_pr__nfet_01v8_lvt_MVT43V
Xsky130_fd_pr__nfet_01v8_lvt_MVT43V_1 m1_964_n363# avss1p8 avss1p8 reg0 avss1p8 sky130_fd_pr__nfet_01v8_lvt_MVT43V
Xsky130_fd_pr__nfet_01v8_lvt_NMSMYT_0 vctrl m1_1996_n363# vctrl avss1p8 m1_1996_n363#
+ iref m1_1996_n363# vctrl m1_1996_n363# vctrl vctrl sky130_fd_pr__nfet_01v8_lvt_NMSMYT
Xsky130_fd_pr__nfet_01v8_lvt_NMSMYT_1 avss1p8 m1_1996_n363# avss1p8 avss1p8 m1_1996_n363#
+ reg2 m1_1996_n363# avss1p8 m1_1996_n363# avss1p8 avss1p8 sky130_fd_pr__nfet_01v8_lvt_NMSMYT
Xsky130_fd_pr__nfet_01v8_lvt_72JNYZ_0 m1_448_n363# avss1p8 iref m1_448_n363# vctrl
+ vctrl sky130_fd_pr__nfet_01v8_lvt_72JNYZ
Xsky130_fd_pr__nfet_01v8_lvt_72JNYZ_1 m1_448_n363# avss1p8 avdd1p8 m1_448_n363# avss1p8
+ avss1p8 sky130_fd_pr__nfet_01v8_lvt_72JNYZ
Xsky130_fd_pr__pfet_01v8_XAYTAL_0 avss1p8 avdd1p8 m1_511_801# avss1p8 m1_511_801#
+ avdd1p8 avdd1p8 sky130_fd_pr__pfet_01v8_XAYTAL
Xsky130_fd_pr__nfet_01v8_lvt_B2JNY3_0 vctrl m1_1384_n363# vctrl m1_1384_n363# avss1p8
+ iref vctrl sky130_fd_pr__nfet_01v8_lvt_B2JNY3
Xsky130_fd_pr__nfet_01v8_lvt_B2JNY3_1 avss1p8 m1_1384_n363# avss1p8 m1_1384_n363#
+ avss1p8 reg1 avss1p8 sky130_fd_pr__nfet_01v8_lvt_B2JNY3
Xsky130_fd_pr__pfet_01v8_XACJHL_0 avss1p8 vctrl avdd1p8 m1_511_801# vctrl vctrl sky130_fd_pr__pfet_01v8_XACJHL
.ends

.subckt res_amp_lin_prog avdd1p8 delay_reg2 clk avss1p8 outp_cap iref_reg0 iref_reg1
+ iref_reg2 iref delay_reg0 inn outn_cap inp delay_reg1 rst
Xsky130_fd_pr__pfet_01v8_lvt_4L9VGG_0 avss1p8 outn_cap avdd1p8 outn_cap res_amp_lin_0/clk
+ outn outn outn outn_cap sky130_fd_pr__pfet_01v8_lvt_4L9VGG
Xsky130_fd_pr__pfet_01v8_lvt_4L9VGG_1 avss1p8 outp_cap avdd1p8 outp_cap res_amp_lin_0/clk
+ outp outp outp outp_cap sky130_fd_pr__pfet_01v8_lvt_4L9VGG
Xdelay_cell_buff_0 clk res_amp_lin_0/clk avss1p8 avdd1p8 delay_reg0 delay_reg2 delay_reg1
+ avss1p8 delay_cell_buff
Xinverter_min_x4_0 avdd1p8 res_amp_lin_0/clk avss1p8 inverter_min_x4_0/out inverter_min_x4
Xsky130_fd_pr__nfet_01v8_lvt_72JNYZ_0 outn_cap avss1p8 rst outn_cap avss1p8 avss1p8
+ sky130_fd_pr__nfet_01v8_lvt_72JNYZ
Xres_amp_lin_0 res_amp_lin_0/clk res_amp_lin_0/vctrl avdd1p8 avss1p8 inn outn outp
+ inp res_amp_lin
Xsky130_fd_pr__nfet_01v8_lvt_72JNYZ_1 outp_cap avss1p8 rst outp_cap avss1p8 avss1p8
+ sky130_fd_pr__nfet_01v8_lvt_72JNYZ
Xsky130_fd_pr__nfet_01v8_lvt_595QY5_0 outn outn outn outn_cap outn_cap avss1p8 outn_cap
+ inverter_min_x4_0/out sky130_fd_pr__nfet_01v8_lvt_595QY5
Xsky130_fd_pr__nfet_01v8_lvt_595QY5_1 outp outp outp outp_cap outp_cap avss1p8 outp_cap
+ inverter_min_x4_0/out sky130_fd_pr__nfet_01v8_lvt_595QY5
Xiref_ctrl_res_amp_0 res_amp_lin_0/vctrl avdd1p8 iref_reg0 iref_reg1 iref_reg2 iref
+ avss1p8 iref_ctrl_res_amp
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_D3F744 VSUBS a_n285_n236# a_355_n236# a_n29_n236#
+ a_n413_n236# a_99_n236# a_n611_n262# a_483_n236# a_n669_n236# w_n807_n384# a_n157_n236#
+ a_n541_n236# a_227_n236# a_611_n236#
X0 a_n157_n236# a_n611_n262# a_n285_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X1 a_611_n236# a_n611_n262# a_483_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X2 a_227_n236# a_n611_n262# a_99_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X3 a_n285_n236# a_n611_n262# a_n413_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X4 a_99_n236# a_n611_n262# a_n29_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X5 a_355_n236# a_n611_n262# a_227_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X6 a_483_n236# a_n611_n262# a_355_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X7 a_n29_n236# a_n611_n262# a_n157_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X8 a_n413_n236# a_n611_n262# a_n541_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
X9 a_n541_n236# a_n611_n262# a_n669_n236# w_n807_n384# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=350000u
.ends

.subckt sky130_fd_pr__pfet_01v8_VCU74W VSUBS a_495_n100# a_n81_n100# a_399_n100# a_687_n100#
+ a_n749_n100# a_n273_n100# a_111_n100# a_n177_n100# a_n561_n100# a_15_n100# a_n465_n100#
+ a_n705_n197# a_303_n100# a_n369_n100# w_n887_n319# a_207_n100# a_n657_n100# a_591_n100#
X0 a_303_n100# a_n705_n197# a_207_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_591_n100# a_n705_n197# a_495_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_207_n100# a_n705_n197# a_111_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_399_n100# a_n705_n197# a_303_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_495_n100# a_n705_n197# a_399_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_687_n100# a_n705_n197# a_591_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n561_n100# a_n705_n197# a_n657_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n465_n100# a_n705_n197# a_n561_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n657_n100# a_n705_n197# a_n749_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n369_n100# a_n705_n197# a_n465_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_15_n100# a_n705_n197# a_n81_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_111_n100# a_n705_n197# a_15_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n273_n100# a_n705_n197# a_n369_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n81_n100# a_n705_n197# a_n177_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n177_n100# a_n705_n197# a_n273_n100# w_n887_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt source_follower_buff_pmos in avdd1p8 out iref avss1p8
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_0 avss1p8 iref iref iref avss1p8 avss1p8 avss1p8
+ avss1p8 iref sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_1 avss1p8 m1_957_828# m1_957_828# iref avss1p8
+ avss1p8 avss1p8 avss1p8 m1_957_828# sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__pfet_01v8_lvt_D3F744_0 avss1p8 out avss1p8 out avss1p8 avss1p8 in out
+ avss1p8 avdd1p8 avss1p8 out out avss1p8 sky130_fd_pr__pfet_01v8_lvt_D3F744
Xsky130_fd_pr__pfet_01v8_VCU74W_0 avss1p8 m1_957_828# m1_957_828# avdd1p8 m1_957_828#
+ avdd1p8 m1_957_828# m1_957_828# avdd1p8 avdd1p8 avdd1p8 m1_957_828# m1_957_828#
+ m1_957_828# avdd1p8 avdd1p8 avdd1p8 m1_957_828# avdd1p8 sky130_fd_pr__pfet_01v8_VCU74W
Xsky130_fd_pr__pfet_01v8_VCU74W_1 avss1p8 out out avdd1p8 out avdd1p8 out out avdd1p8
+ avdd1p8 avdd1p8 out m1_957_828# out avdd1p8 avdd1p8 avdd1p8 out avdd1p8 sky130_fd_pr__pfet_01v8_VCU74W
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_CFLRKA a_n993_109# a_n1473_n309# a_63_n309# a_1215_n309#
+ a_1215_109# a_n129_n309# a_735_109# a_1599_109# a_n513_n309# a_255_109# a_n1377_n309#
+ a_n1949_109# a_n1761_n309# a_1119_n309# a_1503_n309# a_n1761_109# a_n417_109# a_n417_n309#
+ a_n1281_109# a_n801_n309# a_351_n309# a_63_109# a_1503_109# a_n1665_n309# a_1023_109#
+ a_1887_109# a_1407_n309# a_543_109# a_n705_n309# a_255_n309# a_1791_n309# a_n1569_109#
+ a_n705_109# a_n1569_n309# a_n1089_109# w_n2087_n519# a_n225_109# a_n609_n309# a_159_n309#
+ a_543_n309# a_1695_n309# a_1311_109# a_831_109# a_1695_109# a_n1857_n309# a_n993_n309#
+ a_n33_109# a_351_109# a_n1857_109# a_447_n309# a_831_n309# a_1599_n309# a_n1377_109#
+ a_n897_n309# a_n897_109# a_n513_109# a_1119_109# a_639_109# a_n33_n309# a_735_n309#
+ a_1887_n309# a_159_109# a_n1665_109# a_n1281_n309# a_1023_n309# a_n1185_109# a_n801_109#
+ a_639_n309# a_n321_109# a_1407_109# a_n321_n309# a_927_109# a_447_109# a_1791_109#
+ a_n1185_n309# a_1311_n309# a_n1905_n87# a_927_n309# a_n609_109# a_n225_n309# a_n1473_109#
+ a_n129_109# a_n1949_n309# a_n1089_n309#
X0 a_n1569_n309# a_n1905_n87# a_n1665_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n897_n309# a_n1905_n87# a_n993_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_927_n309# a_n1905_n87# a_831_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_1023_109# a_n1905_n87# a_927_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_255_n309# a_n1905_n87# a_159_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1215_n309# a_n1905_n87# a_1119_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_927_109# a_n1905_n87# a_831_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n1857_n309# a_n1905_n87# a_n1949_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n321_n309# a_n1905_n87# a_n417_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n1761_109# a_n1905_n87# a_n1857_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_543_n309# a_n1905_n87# a_447_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_1503_n309# a_n1905_n87# a_1407_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n1857_109# a_n1905_n87# a_n1949_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n1665_109# a_n1905_n87# a_n1761_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n1569_109# a_n1905_n87# a_n1665_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1215_109# a_n1905_n87# a_1119_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_1311_109# a_n1905_n87# a_1215_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_1503_109# a_n1905_n87# a_1407_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_1791_109# a_n1905_n87# a_1695_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n1185_n309# a_n1905_n87# a_n1281_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_1119_109# a_n1905_n87# a_1023_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1407_109# a_n1905_n87# a_1311_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1599_109# a_n1905_n87# a_1503_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_1695_109# a_n1905_n87# a_1599_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_1887_109# a_n1905_n87# a_1791_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_n1473_n309# a_n1905_n87# a_n1569_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_831_n309# a_n1905_n87# a_735_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_1791_n309# a_n1905_n87# a_1695_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n33_109# a_n1905_n87# a_n129_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_351_109# a_n1905_n87# a_255_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_159_n309# a_n1905_n87# a_63_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1119_n309# a_n1905_n87# a_1023_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_159_109# a_n1905_n87# a_63_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_255_109# a_n1905_n87# a_159_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_447_109# a_n1905_n87# a_351_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_543_109# a_n1905_n87# a_447_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_735_109# a_n1905_n87# a_639_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_831_109# a_n1905_n87# a_735_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n225_n309# a_n1905_n87# a_n321_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_639_109# a_n1905_n87# a_543_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_447_n309# a_n1905_n87# a_351_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_1407_n309# a_n1905_n87# a_1311_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_n1473_109# a_n1905_n87# a_n1569_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 a_n1281_109# a_n1905_n87# a_n1377_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 a_n1185_109# a_n1905_n87# a_n1281_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 a_n993_109# a_n1905_n87# a_n1089_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 a_n1089_n309# a_n1905_n87# a_n1185_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 a_n1377_109# a_n1905_n87# a_n1473_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_n1089_109# a_n1905_n87# a_n1185_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 a_n321_109# a_n1905_n87# a_n417_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n513_n309# a_n1905_n87# a_n609_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 a_63_n309# a_n1905_n87# a_n33_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_n801_109# a_n1905_n87# a_n897_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 a_n705_109# a_n1905_n87# a_n801_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_n513_109# a_n1905_n87# a_n609_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_n417_109# a_n1905_n87# a_n513_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 a_n225_109# a_n1905_n87# a_n321_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 a_n129_109# a_n1905_n87# a_n225_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_n1377_n309# a_n1905_n87# a_n1473_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 a_735_n309# a_n1905_n87# a_639_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X60 a_1695_n309# a_n1905_n87# a_1599_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 a_n897_109# a_n1905_n87# a_n993_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 a_n609_109# a_n1905_n87# a_n705_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 a_n801_n309# a_n1905_n87# a_n897_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 a_n129_n309# a_n1905_n87# a_n225_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 a_n1761_n309# a_n1905_n87# a_n1857_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 a_n417_n309# a_n1905_n87# a_n513_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 a_63_109# a_n1905_n87# a_n33_109# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 a_639_n309# a_n1905_n87# a_543_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 a_1599_n309# a_n1905_n87# a_1503_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 a_n705_n309# a_n1905_n87# a_n801_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X71 a_1887_n309# a_n1905_n87# a_1791_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 a_n1665_n309# a_n1905_n87# a_n1761_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 a_1023_n309# a_n1905_n87# a_927_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 a_n993_n309# a_n1905_n87# a_n1089_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 a_n33_n309# a_n1905_n87# a_n129_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 a_351_n309# a_n1905_n87# a_255_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 a_1311_n309# a_n1905_n87# a_1215_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 a_n1281_n309# a_n1905_n87# a_n1377_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X79 a_n609_n309# a_n1905_n87# a_n705_n309# w_n2087_n519# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_CAF2P9 a_63_n309# a_n1473_n309# a_159_527# a_1215_n309#
+ a_n993_109# a_1215_109# a_n129_n309# a_n513_n309# a_1599_109# a_735_109# a_n1665_527#
+ a_n1281_n727# a_n801_527# a_1023_n727# a_639_n727# a_255_109# a_n1185_527# a_n1377_n309#
+ a_n1949_109# a_1119_n309# a_n1761_n309# a_n321_527# a_1503_n309# a_1407_527# a_n321_n727#
+ a_927_527# a_n1761_109# a_n417_109# a_n417_n309# a_351_n309# a_n801_n309# a_n1905_n505#
+ a_n1281_109# a_n1185_n727# a_447_527# a_1791_527# a_63_109# a_1311_n727# a_927_n727#
+ a_1503_109# a_n1665_n309# a_1407_n309# a_1887_109# a_n225_n727# a_1023_109# a_n609_527#
+ a_543_109# a_255_n309# a_n1473_527# a_n1949_n727# a_1791_n309# a_n705_n309# a_n129_527#
+ a_n1089_n727# a_n1473_n727# a_1215_n727# a_63_n727# a_n993_527# a_n1569_109# a_n1569_n309#
+ a_n705_109# a_1215_527# a_n129_n727# a_n1089_109# a_1599_527# a_n513_n727# a_735_527#
+ a_n225_109# a_1695_n309# a_159_n309# a_n609_n309# a_543_n309# a_255_527# a_n1377_n727#
+ a_n1949_527# a_1119_n727# a_n1761_n727# a_1503_n727# a_1311_109# a_n993_n309# a_1695_109#
+ a_n1857_n309# a_831_109# a_n1761_527# a_n33_109# a_n417_n727# a_n417_527# a_351_109#
+ a_351_n727# a_n801_n727# a_n1281_527# a_n1857_109# a_1599_n309# a_447_n309# a_63_527#
+ a_831_n309# a_1503_527# a_n1377_109# a_n1665_n727# a_1887_527# a_1407_n727# a_n897_n309#
+ a_1023_527# a_n513_109# a_n897_109# a_543_527# a_1791_n727# a_255_n727# a_n705_n727#
+ a_1119_109# a_1887_n309# a_639_109# a_735_n309# a_n33_n309# a_n1569_527# a_n1569_n727#
+ a_n705_527# a_159_109# a_n1089_527# a_n225_527# w_n2087_n937# a_1695_n727# a_159_n727#
+ a_n609_n727# a_543_n727# a_n1665_109# a_n1281_n309# a_1023_n309# a_1311_527# a_n801_109#
+ a_639_n309# a_1695_527# a_n1185_109# a_n993_n727# a_831_527# a_n1857_n727# a_n321_109#
+ a_1407_109# a_n33_527# a_n321_n309# a_351_527# a_927_109# a_1599_n727# a_n1857_527#
+ a_447_n727# a_831_n727# a_447_109# a_n1185_n309# a_n1377_527# a_1791_109# a_1311_n309#
+ a_n897_n727# a_927_n309# a_n513_527# a_n897_527# a_n225_n309# a_n609_109# a_1119_527#
+ a_1887_n727# a_n1949_n309# a_639_527# a_n1473_109# a_n129_109# a_735_n727# a_n33_n727#
+ a_n1089_n309#
X0 a_927_n309# a_n1905_n505# a_831_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_n897_n309# a_n1905_n505# a_n993_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n1569_n309# a_n1905_n505# a_n1665_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n129_n727# a_n1905_n505# a_n225_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n1761_n727# a_n1905_n505# a_n1857_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1215_n309# a_n1905_n505# a_1119_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_255_n309# a_n1905_n505# a_159_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_1023_109# a_n1905_n505# a_927_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n1857_n309# a_n1905_n505# a_n1949_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_927_109# a_n1905_n505# a_831_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n417_n727# a_n1905_n505# a_n513_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n321_n309# a_n1905_n505# a_n417_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_1599_n727# a_n1905_n505# a_1503_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_63_527# a_n1905_n505# a_n33_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n1761_109# a_n1905_n505# a_n1857_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1503_n309# a_n1905_n505# a_1407_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_639_n727# a_n1905_n505# a_543_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_543_n309# a_n1905_n505# a_447_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n1665_109# a_n1905_n505# a_n1761_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n1185_n309# a_n1905_n505# a_n1281_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_n1569_109# a_n1905_n505# a_n1665_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1311_109# a_n1905_n505# a_1215_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_n1857_109# a_n1905_n505# a_n1949_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_1791_109# a_n1905_n505# a_1695_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_1503_109# a_n1905_n505# a_1407_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_1215_109# a_n1905_n505# a_1119_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_n705_n727# a_n1905_n505# a_n801_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_1119_109# a_n1905_n505# a_1023_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1695_109# a_n1905_n505# a_1599_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1407_109# a_n1905_n505# a_1311_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_1599_109# a_n1905_n505# a_1503_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1887_109# a_n1905_n505# a_1791_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1887_n727# a_n1905_n505# a_1791_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_1791_n309# a_n1905_n505# a_1695_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_831_n309# a_n1905_n505# a_735_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_n1473_n309# a_n1905_n505# a_n1569_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_n33_109# a_n1905_n505# a_n129_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_1023_n727# a_n1905_n505# a_927_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n1665_n727# a_n1905_n505# a_n1761_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_1119_n309# a_n1905_n505# a_1023_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_159_n309# a_n1905_n505# a_63_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_351_109# a_n1905_n505# a_255_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_1311_n727# a_n1905_n505# a_1215_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 a_255_109# a_n1905_n505# a_159_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 a_351_n727# a_n1905_n505# a_255_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 a_831_109# a_n1905_n505# a_735_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 a_543_109# a_n1905_n505# a_447_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 a_n33_n727# a_n1905_n505# a_n129_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_n993_n727# a_n1905_n505# a_n1089_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 a_159_109# a_n1905_n505# a_63_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n225_n309# a_n1905_n505# a_n321_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 a_735_109# a_n1905_n505# a_639_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_447_109# a_n1905_n505# a_351_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 a_639_109# a_n1905_n505# a_543_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_1407_n309# a_n1905_n505# a_1311_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_447_n309# a_n1905_n505# a_351_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 a_n1089_n309# a_n1905_n505# a_n1185_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 a_n1281_109# a_n1905_n505# a_n1377_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_n993_109# a_n1905_n505# a_n1089_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 a_n1473_109# a_n1905_n505# a_n1569_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X60 a_n1185_109# a_n1905_n505# a_n1281_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 a_n609_n727# a_n1905_n505# a_n705_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 a_n1377_109# a_n1905_n505# a_n1473_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 a_n1089_109# a_n1905_n505# a_n1185_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 a_n1281_n727# a_n1905_n505# a_n1377_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 a_n513_n309# a_n1905_n505# a_n609_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 a_n321_109# a_n1905_n505# a_n417_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 a_63_n309# a_n1905_n505# a_n33_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 a_n225_109# a_n1905_n505# a_n321_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 a_n801_109# a_n1905_n505# a_n897_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 a_n513_109# a_n1905_n505# a_n609_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X71 a_1695_n309# a_n1905_n505# a_1599_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 a_n705_109# a_n1905_n505# a_n801_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 a_n417_109# a_n1905_n505# a_n513_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 a_n129_109# a_n1905_n505# a_n225_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 a_735_n309# a_n1905_n505# a_639_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 a_n1377_n309# a_n1905_n505# a_n1473_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 a_n897_109# a_n1905_n505# a_n993_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 a_n609_109# a_n1905_n505# a_n705_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X79 a_927_n727# a_n1905_n505# a_831_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X80 a_n1569_n727# a_n1905_n505# a_n1665_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X81 a_n897_n727# a_n1905_n505# a_n993_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X82 a_n801_n309# a_n1905_n505# a_n897_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 a_1215_n727# a_n1905_n505# a_1119_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X84 a_255_n727# a_n1905_n505# a_159_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X85 a_1023_527# a_n1905_n505# a_927_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X86 a_n129_n309# a_n1905_n505# a_n225_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X87 a_927_527# a_n1905_n505# a_831_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X88 a_n1857_n727# a_n1905_n505# a_n1949_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X89 a_n1761_n309# a_n1905_n505# a_n1857_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X90 a_n321_n727# a_n1905_n505# a_n417_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X91 a_n1761_527# a_n1905_n505# a_n1857_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 a_1503_n727# a_n1905_n505# a_1407_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X93 a_n1665_527# a_n1905_n505# a_n1761_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X94 a_543_n727# a_n1905_n505# a_447_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X95 a_n1185_n727# a_n1905_n505# a_n1281_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X96 a_n417_n309# a_n1905_n505# a_n513_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X97 a_n1857_527# a_n1905_n505# a_n1949_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X98 a_n1569_527# a_n1905_n505# a_n1665_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 a_1311_527# a_n1905_n505# a_1215_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X100 a_1215_527# a_n1905_n505# a_1119_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 a_1503_527# a_n1905_n505# a_1407_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X102 a_1791_527# a_n1905_n505# a_1695_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X103 a_1119_527# a_n1905_n505# a_1023_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X104 a_1407_527# a_n1905_n505# a_1311_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X105 a_1695_527# a_n1905_n505# a_1599_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X106 a_1599_n309# a_n1905_n505# a_1503_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X107 a_63_109# a_n1905_n505# a_n33_109# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X108 a_639_n309# a_n1905_n505# a_543_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X109 a_1599_527# a_n1905_n505# a_1503_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X110 a_1887_527# a_n1905_n505# a_1791_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X111 a_1791_n727# a_n1905_n505# a_1695_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X112 a_831_n727# a_n1905_n505# a_735_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X113 a_n1473_n727# a_n1905_n505# a_n1569_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 a_n705_n309# a_n1905_n505# a_n801_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 a_n33_527# a_n1905_n505# a_n129_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 a_1887_n309# a_n1905_n505# a_1791_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X117 a_1119_n727# a_n1905_n505# a_1023_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 a_159_n727# a_n1905_n505# a_63_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X119 a_351_527# a_n1905_n505# a_255_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X120 a_1023_n309# a_n1905_n505# a_927_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X121 a_n1665_n309# a_n1905_n505# a_n1761_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X122 a_255_527# a_n1905_n505# a_159_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X123 a_543_527# a_n1905_n505# a_447_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X124 a_831_527# a_n1905_n505# a_735_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X125 a_159_527# a_n1905_n505# a_63_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X126 a_447_527# a_n1905_n505# a_351_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X127 a_n225_n727# a_n1905_n505# a_n321_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X128 a_735_527# a_n1905_n505# a_639_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X129 a_639_527# a_n1905_n505# a_543_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X130 a_1407_n727# a_n1905_n505# a_1311_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X131 a_447_n727# a_n1905_n505# a_351_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X132 a_1311_n309# a_n1905_n505# a_1215_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X133 a_n1089_n727# a_n1905_n505# a_n1185_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X134 a_351_n309# a_n1905_n505# a_255_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 a_n33_n309# a_n1905_n505# a_n129_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X136 a_n1281_527# a_n1905_n505# a_n1377_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X137 a_n993_527# a_n1905_n505# a_n1089_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X138 a_n993_n309# a_n1905_n505# a_n1089_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X139 a_n1473_527# a_n1905_n505# a_n1569_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 a_n1185_527# a_n1905_n505# a_n1281_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X141 a_n1377_527# a_n1905_n505# a_n1473_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X142 a_n1089_527# a_n1905_n505# a_n1185_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X143 a_n513_n727# a_n1905_n505# a_n609_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X144 a_n321_527# a_n1905_n505# a_n417_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X145 a_63_n727# a_n1905_n505# a_n33_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X146 a_n801_527# a_n1905_n505# a_n897_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X147 a_n513_527# a_n1905_n505# a_n609_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X148 a_n225_527# a_n1905_n505# a_n321_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X149 a_1695_n727# a_n1905_n505# a_1599_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X150 a_735_n727# a_n1905_n505# a_639_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X151 a_n705_527# a_n1905_n505# a_n801_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X152 a_n417_527# a_n1905_n505# a_n513_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X153 a_n129_527# a_n1905_n505# a_n225_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X154 a_n1377_n727# a_n1905_n505# a_n1473_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 a_n609_n309# a_n1905_n505# a_n705_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 a_n1281_n309# a_n1905_n505# a_n1377_n309# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X157 a_n897_527# a_n1905_n505# a_n993_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X158 a_n609_527# a_n1905_n505# a_n705_527# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X159 a_n801_n727# a_n1905_n505# a_n897_n727# w_n2087_n937# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt source_follower_buff_nmos in avdd1p8 avss1p8 out iref
Xsky130_fd_pr__nfet_01v8_lvt_CFLRKA_0 avdd1p8 out out out out out avdd1p8 out out
+ out avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 out avdd1p8
+ avdd1p8 out avdd1p8 out out avdd1p8 out avdd1p8 out out out avdd1p8 out avdd1p8
+ out avss1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 avdd1p8 out avdd1p8 out avdd1p8
+ avdd1p8 avdd1p8 out out out out avdd1p8 out out out avdd1p8 out avdd1p8 avdd1p8
+ avdd1p8 avdd1p8 out out out avdd1p8 avdd1p8 out out out out avdd1p8 out out avdd1p8
+ avdd1p8 in avdd1p8 avdd1p8 avdd1p8 out out avdd1p8 out sky130_fd_pr__nfet_01v8_lvt_CFLRKA
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_0 m1_460_n1129# iref iref iref m1_460_n1129# m1_460_n1129#
+ avss1p8 m1_460_n1129# iref sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_9B2JY7_1 avss1p8 m1_460_n1129# m1_460_n1129# iref avss1p8
+ avss1p8 avss1p8 avss1p8 m1_460_n1129# sky130_fd_pr__nfet_01v8_lvt_9B2JY7
Xsky130_fd_pr__nfet_01v8_lvt_CAF2P9_0 out out avss1p8 out avss1p8 out out out out
+ avss1p8 out out avss1p8 out out out avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 out
+ avss1p8 out out avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 iref out avss1p8
+ out out out avss1p8 avss1p8 avss1p8 out out avss1p8 avss1p8 out avss1p8 avss1p8
+ out out avss1p8 out out out out out out out avss1p8 avss1p8 avss1p8 out out out
+ out out out avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 out avss1p8 avss1p8
+ avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 out out avss1p8 avss1p8 avss1p8
+ avss1p8 avss1p8 avss1p8 avss1p8 out out out out out out avss1p8 avss1p8 out avss1p8
+ out out out out out avss1p8 out out out avss1p8 avss1p8 out avss1p8 avss1p8 avss1p8
+ avss1p8 out avss1p8 out avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 avss1p8 out out
+ out avss1p8 avss1p8 out avss1p8 avss1p8 avss1p8 out out out out avss1p8 out avss1p8
+ avss1p8 out out out out out avss1p8 avss1p8 out avss1p8 out avss1p8 out out avss1p8
+ avss1p8 avss1p8 avss1p8 avss1p8 out out out avss1p8 avss1p8 out sky130_fd_pr__nfet_01v8_lvt_CAF2P9
.ends

.subckt source_follower_buff_diff VSUBS avdd1p8 iref1 iref2 iref3 iref4 inn outn inp
+ outp
Xsource_follower_buff_pmos_0 inn avdd1p8 source_follower_buff_nmos_0/in iref3 VSUBS
+ source_follower_buff_pmos
Xsource_follower_buff_pmos_1 inp avdd1p8 source_follower_buff_nmos_1/in iref1 VSUBS
+ source_follower_buff_pmos
Xsource_follower_buff_nmos_0 source_follower_buff_nmos_0/in avdd1p8 VSUBS outn iref4
+ source_follower_buff_nmos
Xsource_follower_buff_nmos_1 source_follower_buff_nmos_1/in avdd1p8 VSUBS outp iref2
+ source_follower_buff_nmos
.ends

.subckt res_amp_top iref0 iref1 avss1p8 iref2 iref3 iref4 avdd1p8 res_amp_sync_v2_0/clkp
+ iref_reg0 iref_reg1 iref_reg2 delay_reg0 delay_reg1 inn outn delay_reg2 outp inp
+ clkn
Xres_amp_sync_v2_0 avss1p8 avdd1p8 res_amp_lin_prog_0/clk clkn res_amp_sync_v2_0/clkp
+ res_amp_sync_v2_0/rst res_amp_sync_v2
Xres_amp_lin_prog_0 avdd1p8 delay_reg2 res_amp_lin_prog_0/clk avss1p8 res_amp_lin_prog_0/outp_cap
+ iref_reg0 iref_reg1 iref_reg2 iref0 delay_reg0 inn res_amp_lin_prog_0/outn_cap inp
+ delay_reg1 res_amp_sync_v2_0/rst res_amp_lin_prog
Xsource_follower_buff_diff_0 avss1p8 avdd1p8 iref1 iref2 iref3 iref4 res_amp_lin_prog_0/outn_cap
+ outn res_amp_lin_prog_0/outp_cap outp source_follower_buff_diff
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MACBVW VSUBS m3_n2650_n13200# m3_n7969_n2600# m3_7988_8000#
+ m3_2669_n7900# m3_n13288_n2600# m3_n2650_2700# m3_2669_2700# m3_n13288_n13200# m3_n7969_n13200#
+ m3_n13288_8000# m3_7988_2700# m3_n2650_n7900# m3_7988_n7900# m3_2669_n13200# m3_n7969_8000#
+ m3_n13288_2700# m3_n7969_n7900# m3_n13288_n7900# m3_2669_n2600# m3_n7969_2700# m3_7988_n13200#
+ c1_n13188_n13100# m3_7988_n2600# m3_n2650_n2600# m3_n2650_8000# m3_2669_8000#
X0 c1_n13188_n13100# m3_2669_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X1 c1_n13188_n13100# m3_n2650_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X2 c1_n13188_n13100# m3_2669_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X3 c1_n13188_n13100# m3_n13288_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X4 c1_n13188_n13100# m3_n7969_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X5 c1_n13188_n13100# m3_n13288_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X6 c1_n13188_n13100# m3_2669_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X7 c1_n13188_n13100# m3_7988_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X8 c1_n13188_n13100# m3_2669_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X9 c1_n13188_n13100# m3_7988_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X10 c1_n13188_n13100# m3_n7969_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X11 c1_n13188_n13100# m3_7988_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X12 c1_n13188_n13100# m3_n7969_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X13 c1_n13188_n13100# m3_7988_8000# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X14 c1_n13188_n13100# m3_n13288_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X15 c1_n13188_n13100# m3_n7969_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X16 c1_n13188_n13100# m3_n2650_n7900# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X17 c1_n13188_n13100# m3_n2650_n13200# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X18 c1_n13188_n13100# m3_n2650_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X19 c1_n13188_n13100# m3_7988_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X20 c1_n13188_n13100# m3_n13288_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X21 c1_n13188_n13100# m3_n13288_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X22 c1_n13188_n13100# m3_n7969_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X23 c1_n13188_n13100# m3_n2650_n2600# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X24 c1_n13188_n13100# m3_2669_2700# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
.ends

.subckt cap1_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_MACBVW_0 VSUBS out out out out out out out out out out
+ out out out out out out out out out out out in out out out out sky130_fd_pr__cap_mim_m3_1_MACBVW
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_W3JTNJ VSUBS m3_n6469_n2100# c1_n6369_n6300# m3_2169_n6400#
+ m3_n2150_n6400# c1_2269_n6300# m3_n6469_2200# m3_n2150_n2100# c1_n2050_n6300# m3_n2150_2200#
+ m3_n6469_n6400#
X0 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2 c1_n2050_n6300# m3_n2150_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 c1_n6369_n6300# m3_n6469_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X4 c1_2269_n6300# m3_2169_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X5 c1_n6369_n6300# m3_n6469_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X6 c1_n2050_n6300# m3_n2150_n2100# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X7 c1_n2050_n6300# m3_n2150_n6400# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X8 c1_n6369_n6300# m3_n6469_2200# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
.ends

.subckt cap2_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_W3JTNJ_0 VSUBS out in out out in out out in out out sky130_fd_pr__cap_mim_m3_1_W3JTNJ
.ends

.subckt sky130_fd_pr__res_high_po_5p73_X44RQA a_n573_2292# w_n739_n2890# a_n573_n2724#
X0 a_n573_n2724# a_n573_2292# w_n739_n2890# sky130_fd_pr__res_high_po_5p73 l=2.292e+07u
.ends

.subckt res_loop_filter vss out in
Xsky130_fd_pr__res_high_po_5p73_X44RQA_0 in vss out sky130_fd_pr__res_high_po_5p73_X44RQA
.ends

.subckt loop_filter vc_pex in vss
Xcap1_loop_filter_0 vss vc_pex vss cap1_loop_filter
Xcap2_loop_filter_0 vss in vss cap2_loop_filter
Xres_loop_filter_0 vss res_loop_filter_2/out in res_loop_filter
Xres_loop_filter_1 vss res_loop_filter_2/out vc_pex res_loop_filter
Xres_loop_filter_2 vss res_loop_filter_2/out vc_pex res_loop_filter
.ends

.subckt sky130_fd_pr__pfet_01v8_4ML9WA VSUBS a_429_n486# w_n2457_n634# a_887_n486#
+ a_n29_n486# a_1345_n486# a_n2261_n512# a_1803_n486# a_n487_n486# a_n945_n486# a_n2319_n486#
+ a_n1403_n486# a_2261_n486# a_n1861_n486#
X0 a_2261_n486# a_n2261_n512# a_1803_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X1 a_n945_n486# a_n2261_n512# a_n1403_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X2 a_429_n486# a_n2261_n512# a_n29_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X3 a_1803_n486# a_n2261_n512# a_1345_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X4 a_887_n486# a_n2261_n512# a_429_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X5 a_n487_n486# a_n2261_n512# a_n945_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X6 a_n1403_n486# a_n2261_n512# a_n1861_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X7 a_n1861_n486# a_n2261_n512# a_n2319_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X8 a_n29_n486# a_n2261_n512# a_n487_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
X9 a_1345_n486# a_n2261_n512# a_887_n486# w_n2457_n634# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_YCGG98 a_n1041_n75# a_n561_n75# a_1167_n75# a_303_n75#
+ a_687_n75# a_n849_n75# a_n369_n75# a_975_n75# a_111_n75# a_495_n75# a_n1137_n75#
+ a_n657_n75# a_n177_n75# a_783_n75# a_n945_n75# a_n465_n75# a_207_n75# a_1071_n75#
+ a_591_n75# a_15_n75# a_n753_n75# w_n1367_n285# a_n273_n75# a_879_n75# a_399_n75#
+ a_n1229_n75# a_n81_n75# a_n1167_n101#
X0 a_207_n75# a_n1167_n101# a_111_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_303_n75# a_n1167_n101# a_207_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_399_n75# a_n1167_n101# a_303_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_495_n75# a_n1167_n101# a_399_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_591_n75# a_n1167_n101# a_495_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_783_n75# a_n1167_n101# a_687_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_687_n75# a_n1167_n101# a_591_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_879_n75# a_n1167_n101# a_783_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_975_n75# a_n1167_n101# a_879_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_n1041_n75# a_n1167_n101# a_n1137_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_n1137_n75# a_n1167_n101# a_n1229_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n561_n75# a_n1167_n101# a_n657_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_1071_n75# a_n1167_n101# a_975_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n945_n75# a_n1167_n101# a_n1041_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n753_n75# a_n1167_n101# a_n849_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n657_n75# a_n1167_n101# a_n753_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n465_n75# a_n1167_n101# a_n561_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n369_n75# a_n1167_n101# a_n465_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_1167_n75# a_n1167_n101# a_1071_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n849_n75# a_n1167_n101# a_n945_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X20 a_15_n75# a_n1167_n101# a_n81_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X21 a_n81_n75# a_n1167_n101# a_n177_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X22 a_111_n75# a_n1167_n101# a_15_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X23 a_n273_n75# a_n1167_n101# a_n369_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X24 a_n177_n75# a_n1167_n101# a_n273_n75# w_n1367_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_MUHGM9 a_33_n101# a_n129_n75# a_735_n75# a_255_n75#
+ a_n417_n75# a_n989_n75# a_63_n75# a_543_n75# a_n705_n75# a_n225_n75# a_n33_n75#
+ a_831_n75# a_351_n75# a_n927_n101# a_n513_n75# a_n897_n75# w_n1127_n285# a_639_n75#
+ a_159_n75# a_n801_n75# a_n321_n75# a_927_n75# a_447_n75# a_n609_n75#
X0 a_63_n75# a_33_n101# a_n33_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1 a_927_n75# a_33_n101# a_831_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2 a_n33_n75# a_n927_n101# a_n129_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X3 a_159_n75# a_33_n101# a_63_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_255_n75# a_33_n101# a_159_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X5 a_351_n75# a_33_n101# a_255_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X6 a_447_n75# a_33_n101# a_351_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X7 a_543_n75# a_33_n101# a_447_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X8 a_735_n75# a_33_n101# a_639_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_831_n75# a_33_n101# a_735_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X10 a_639_n75# a_33_n101# a_543_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_n321_n75# a_n927_n101# a_n417_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_n801_n75# a_n927_n101# a_n897_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_n705_n75# a_n927_n101# a_n801_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_n513_n75# a_n927_n101# a_n609_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_n417_n75# a_n927_n101# a_n513_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X16 a_n225_n75# a_n927_n101# a_n321_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X17 a_n129_n75# a_n927_n101# a_n225_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X18 a_n897_n75# a_n927_n101# a_n989_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X19 a_n609_n75# a_n927_n101# a_n705_n75# w_n1127_n285# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_NKZXKB VSUBS a_33_n247# a_n801_n150# a_n417_n150#
+ a_351_n150# a_255_n150# a_n705_n150# a_n609_n150# a_159_n150# a_543_n150# a_447_n150#
+ a_831_n150# a_n897_n150# a_n33_n150# a_735_n150# a_n927_n247# a_639_n150# a_n321_n150#
+ a_927_n150# a_n225_n150# a_63_n150# a_n989_n150# a_n513_n150# a_n129_n150# w_n1127_n369#
X0 a_n513_n150# a_n927_n247# a_n609_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_63_n150# a_33_n247# a_n33_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_735_n150# a_33_n247# a_639_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n801_n150# a_n927_n247# a_n897_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n927_n247# a_n225_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n927_n247# a_n513_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_639_n150# a_33_n247# a_543_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n705_n150# a_n927_n247# a_n801_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n33_n150# a_n927_n247# a_n129_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_351_n150# a_33_n247# a_255_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_n609_n150# a_n927_n247# a_n705_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n897_n150# a_n927_n247# a_n989_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_927_n150# a_33_n247# a_831_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_255_n150# a_33_n247# a_159_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n321_n150# a_n927_n247# a_n417_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_543_n150# a_33_n247# a_447_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_831_n150# a_33_n247# a_735_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_159_n150# a_33_n247# a_63_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_n225_n150# a_n927_n247# a_n321_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_447_n150# a_33_n247# a_351_n150# w_n1127_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_8GRULZ a_n1761_n132# a_1045_n44# a_n1461_n44# a_n1103_n44#
+ a_n29_n44# a_n387_n44# a_1761_n44# a_n1819_n44# a_1403_n44# a_687_n44# w_n1957_n254#
+ a_329_n44# a_n745_n44#
X0 a_329_n44# a_n1761_n132# a_n29_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X1 a_1761_n44# a_n1761_n132# a_1403_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X2 a_n745_n44# a_n1761_n132# a_n1103_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X3 a_1045_n44# a_n1761_n132# a_687_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X4 a_n29_n44# a_n1761_n132# a_n387_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X5 a_n1103_n44# a_n1761_n132# a_n1461_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X6 a_n387_n44# a_n1761_n132# a_n745_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X7 a_687_n44# a_n1761_n132# a_329_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X8 a_1403_n44# a_n1761_n132# a_1045_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
X9 a_n1461_n44# a_n1761_n132# a_n1819_n44# w_n1957_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=1.5e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_ND88ZC VSUBS a_303_n150# a_n753_n150# a_n369_n150#
+ w_n1367_n369# a_207_n150# a_n657_n150# a_591_n150# a_n1229_n150# a_n945_n150# a_495_n150#
+ a_n1041_n150# a_n849_n150# a_n81_n150# a_399_n150# a_783_n150# a_1071_n150# a_687_n150#
+ a_975_n150# a_n1137_n150# a_n273_n150# a_111_n150# a_879_n150# a_n177_n150# a_n561_n150#
+ a_15_n150# a_1167_n150# a_n1167_n247# a_n465_n150#
X0 a_n1137_n150# a_n1167_n247# a_n1229_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_495_n150# a_n1167_n247# a_399_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n561_n150# a_n1167_n247# a_n657_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_111_n150# a_n1167_n247# a_15_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_783_n150# a_n1167_n247# a_687_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_1071_n150# a_n1167_n247# a_975_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_399_n150# a_n1167_n247# a_303_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_n465_n150# a_n1167_n247# a_n561_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_687_n150# a_n1167_n247# a_591_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n753_n150# a_n1167_n247# a_n849_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X10 a_975_n150# a_n1167_n247# a_879_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_n81_n150# a_n1167_n247# a_n177_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_15_n150# a_n1167_n247# a_n81_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_n1041_n150# a_n1167_n247# a_n1137_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 a_n369_n150# a_n1167_n247# a_n465_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 a_n657_n150# a_n1167_n247# a_n753_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X16 a_879_n150# a_n1167_n247# a_783_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X17 a_n945_n150# a_n1167_n247# a_n1041_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X18 a_1167_n150# a_n1167_n247# a_1071_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X19 a_303_n150# a_n1167_n247# a_207_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X20 a_n273_n150# a_n1167_n247# a_n369_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X21 a_591_n150# a_n1167_n247# a_495_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X22 a_n849_n150# a_n1167_n247# a_n945_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X23 a_207_n150# a_n1167_n247# a_111_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X24 a_n177_n150# a_n1167_n247# a_n273_n150# w_n1367_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt charge_pump Down out iref pswitch nDown biasp Up nswitch vss vdd nUp
Xsky130_fd_pr__pfet_01v8_4ML9WA_0 vss pswitch vdd pswitch pswitch pswitch nUp pswitch
+ pswitch pswitch pswitch pswitch pswitch pswitch sky130_fd_pr__pfet_01v8_4ML9WA
Xsky130_fd_pr__nfet_01v8_YCGG98_0 vss out out vss vss vss out out vss vss out vss
+ out out out vss out vss out out out vss vss vss out vss vss nswitch sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_1 iref vss vss iref iref iref vss vss iref iref vss
+ iref vss vss vss iref vss iref vss vss vss vss iref iref vss iref iref iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_YCGG98_2 biasp vss vss biasp biasp biasp vss vss biasp biasp
+ vss biasp vss vss vss biasp vss biasp vss vss vss vss biasp biasp vss biasp biasp
+ iref sky130_fd_pr__nfet_01v8_YCGG98
Xsky130_fd_pr__nfet_01v8_MUHGM9_0 nDown iref nswitch vss nswitch nswitch vss nswitch
+ iref nswitch nswitch vss nswitch Down iref iref vss vss nswitch nswitch iref nswitch
+ vss nswitch sky130_fd_pr__nfet_01v8_MUHGM9
Xsky130_fd_pr__pfet_01v8_NKZXKB_0 vss Up pswitch pswitch pswitch vdd biasp pswitch
+ pswitch pswitch vdd vdd biasp pswitch pswitch nUp vdd biasp pswitch pswitch vdd
+ pswitch biasp biasp vdd sky130_fd_pr__pfet_01v8_NKZXKB
Xsky130_fd_pr__nfet_01v8_8GRULZ_0 Down nswitch nswitch nswitch nswitch nswitch nswitch
+ nswitch nswitch nswitch vss nswitch nswitch sky130_fd_pr__nfet_01v8_8GRULZ
Xsky130_fd_pr__pfet_01v8_ND88ZC_0 vss vdd out out vdd out vdd out vdd out vdd vdd
+ vdd vdd out out vdd vdd out out vdd vdd vdd out out out out pswitch vdd sky130_fd_pr__pfet_01v8_ND88ZC
Xsky130_fd_pr__pfet_01v8_ND88ZC_1 vss biasp vdd vdd vdd vdd biasp vdd biasp vdd biasp
+ biasp biasp biasp vdd vdd biasp biasp vdd vdd biasp biasp biasp vdd vdd vdd vdd
+ biasp biasp sky130_fd_pr__pfet_01v8_ND88ZC
.ends

.subckt sky130_fd_pr__nfet_01v8_5RJ8EK a_n33_n42# a_33_n68# w_n263_n252# a_n63_n68#
+ a_n125_n42# a_63_n42#
X0 a_63_n42# a_33_n68# a_n33_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_n33_n42# a_n63_n68# a_n125_n42# w_n263_n252# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_ZPB9BB VSUBS a_n63_n110# a_33_n110# a_n125_n84# a_63_n84#
+ w_n263_n303# a_n33_n84#
X0 a_63_n84# a_33_n110# a_n33_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_n33_n84# a_n63_n110# a_n125_n84# w_n263_n303# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt inverter_min_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_5RJ8EK_0 vss in vss in out out sky130_fd_pr__nfet_01v8_5RJ8EK
Xsky130_fd_pr__pfet_01v8_ZPB9BB_0 vss in in out out vdd vdd sky130_fd_pr__pfet_01v8_ZPB9BB
.ends

.subckt div_by_2 vss vdd CLK_2 nCLK_2 o1 CLK out_div o2 nout_div
XDFlipFlop_0 vss nout_div out_div nout_div vdd DFlipFlop_0/CLK DFlipFlop_0/nCLK DFlipFlop
Xinverter_min_x4_1 vdd o2 vss nCLK_2 inverter_min_x4
Xinverter_min_x4_0 vdd o1 vss CLK_2 inverter_min_x4
Xclock_inverter_0 vss CLK vdd DFlipFlop_0/CLK DFlipFlop_0/nCLK clock_inverter
Xinverter_min_x2_0 nout_div o2 vss vdd inverter_min_x2
Xinverter_min_x2_1 out_div o1 vss vdd inverter_min_x2
.ends

.subckt sky130_fd_pr__pfet_01v8_58ZKDE VSUBS a_n257_n777# a_n129_n600# a_n221_n600#
+ w_n257_n702#
X0 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X1 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X2 a_n129_n600# a_n257_n777# a_n221_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X3 a_n221_n600# a_n257_n777# a_n129_n600# w_n257_n702# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_T69Y3A a_n129_n300# a_n221_n300# w_n257_n327# a_n257_n404#
X0 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2 a_n129_n300# a_n257_n404# a_n221_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 a_n221_n300# a_n257_n404# a_n129_n300# w_n257_n327# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends

.subckt buffer_salida in out vss vdd
Xsky130_fd_pr__pfet_01v8_58ZKDE_1 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_2 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_3 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_0 a_678_n100# vss vss in sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_1 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_4 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_5 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_2 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_3 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_6 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_70 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_4 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_7 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_8 vss a_678_n100# a_3996_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_71 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_60 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_5 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_72 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_61 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_50 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_6 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_9 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_62 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_51 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_7 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_40 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_8 a_3996_n100# vss vss a_678_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_63 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_52 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_30 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_41 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_64 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_53 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_9 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_20 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_31 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_42 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_65 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_54 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_10 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_21 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_32 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_43 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_66 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_55 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_11 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_22 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_33 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_44 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_67 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_56 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_12 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_23 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_34 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_45 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_68 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_57 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_13 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_24 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_35 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_46 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_69 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_58 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_14 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_25 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_36 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_47 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_59 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_48 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_15 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_26 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_37 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_49 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_16 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_27 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_38 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_70 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_17 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_28 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_39 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_71 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_60 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_18 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__nfet_01v8_T69Y3A_29 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_72 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_61 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_50 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_62 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_51 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__nfet_01v8_T69Y3A_19 out vss vss a_3996_n100# sky130_fd_pr__nfet_01v8_T69Y3A
Xsky130_fd_pr__pfet_01v8_58ZKDE_40 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_63 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_52 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_30 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_41 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_64 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_53 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_20 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_31 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_42 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_65 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_54 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_10 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_21 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_32 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_43 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_66 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_55 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_11 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_22 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_33 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_44 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_67 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_56 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_12 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_23 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_34 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_45 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_68 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_57 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_46 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_13 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_24 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_35 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_69 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_58 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_14 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_25 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_36 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_47 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_59 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_15 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_26 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_37 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_48 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_49 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_16 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_27 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_38 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_17 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_28 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_39 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_18 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_29 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_19 vss a_3996_n100# out vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
Xsky130_fd_pr__pfet_01v8_58ZKDE_0 vss in a_678_n100# vdd vdd sky130_fd_pr__pfet_01v8_58ZKDE
.ends

.subckt sky130_fd_pr__nfet_01v8_CBAU6Y a_n73_n150# a_n33_n238# w_n211_n360# a_15_n150#
X0 a_15_n150# a_n33_n238# a_n73_n150# w_n211_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4757AC VSUBS a_n73_n150# a_n33_181# w_n211_n369# a_15_n150#
X0 a_15_n150# a_n33_181# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_7H8F5S a_n465_172# a_n417_n150# a_351_n150# a_255_n150#
+ w_n647_n360# a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150#
X0 a_159_n150# a_n465_172# a_63_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n225_n150# a_n465_172# a_n321_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_447_n150# a_n465_172# a_351_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_63_n150# a_n465_172# a_n33_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_n129_n150# a_n465_172# a_n225_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n417_n150# a_n465_172# a_n509_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n33_n150# a_n465_172# a_n129_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_351_n150# a_n465_172# a_255_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_255_n150# a_n465_172# a_159_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n321_n150# a_n465_172# a_n417_n150# w_n647_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_8DL6ZL VSUBS a_n417_n150# a_351_n150# a_255_n150#
+ a_159_n150# a_447_n150# a_n509_n150# a_n33_n150# a_n465_n247# a_n321_n150# a_n225_n150#
+ a_63_n150# a_n129_n150# w_n647_n369#
X0 a_63_n150# a_n465_n247# a_n33_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X1 a_n129_n150# a_n465_n247# a_n225_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X2 a_n417_n150# a_n465_n247# a_n509_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X3 a_n33_n150# a_n465_n247# a_n129_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X4 a_351_n150# a_n465_n247# a_255_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_255_n150# a_n465_n247# a_159_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X6 a_n321_n150# a_n465_n247# a_n417_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X7 a_159_n150# a_n465_n247# a_63_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_n225_n150# a_n465_n247# a_n321_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_447_n150# a_n465_n247# a_351_n150# w_n647_n369# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_EDT3AT a_15_n11# a_n33_n99# w_n211_n221# a_n73_n11#
X0 a_15_n11# a_n33_n99# a_n73_n11# w_n211_n221# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_AQR2CW a_n33_66# a_n78_n106# w_n216_n254# a_20_n106#
X0 a_20_n106# a_n33_66# a_n78_n106# w_n216_n254# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=750000u l=200000u
.ends

.subckt sky130_fd_pr__pfet_01v8_HRYSXS VSUBS a_n33_n211# a_n78_n114# w_n216_n334#
+ a_20_n114#
X0 a_20_n114# a_n33_n211# a_n78_n114# w_n216_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=200000u
.ends

.subckt inverter_csvco in vbulkn out vbulkp vdd vss
Xsky130_fd_pr__nfet_01v8_AQR2CW_0 in vss vbulkn out sky130_fd_pr__nfet_01v8_AQR2CW
Xsky130_fd_pr__pfet_01v8_HRYSXS_0 vbulkn in vdd vbulkp out sky130_fd_pr__pfet_01v8_HRYSXS
.ends

.subckt cap_vco t b VSUBS
C0 t b 5.78fF
*C1 t VSUBS 0.42fF
*C2 b VSUBS 0.09fF
.ends


.subckt csvco_branch vctrl in vbp D0 out vss vdd
Xsky130_fd_pr__nfet_01v8_7H8F5S_0 vctrl inverter_csvco_0/vss inverter_csvco_0/vss
+ vss vss inverter_csvco_0/vss vss vss inverter_csvco_0/vss vss inverter_csvco_0/vss
+ vss vss sky130_fd_pr__nfet_01v8_7H8F5S
Xsky130_fd_pr__pfet_01v8_8DL6ZL_0 vss inverter_csvco_0/vdd inverter_csvco_0/vdd vdd
+ inverter_csvco_0/vdd vdd vdd inverter_csvco_0/vdd vbp vdd inverter_csvco_0/vdd vdd
+ vdd vdd sky130_fd_pr__pfet_01v8_8DL6ZL
Xsky130_fd_pr__nfet_01v8_EDT3AT_0 cap_vco_0/t D0 vss out sky130_fd_pr__nfet_01v8_EDT3AT
Xinverter_csvco_0 in vss out vdd inverter_csvco_0/vdd inverter_csvco_0/vss inverter_csvco
Xcap_vco_0 cap_vco_0/t vss vss cap_vco
.ends

.subckt ring_osc vctrl vdd vss D0 out_vco
Xsky130_fd_pr__nfet_01v8_CBAU6Y_0 vss vctrl vss csvco_branch_2/vbp sky130_fd_pr__nfet_01v8_CBAU6Y
Xsky130_fd_pr__pfet_01v8_4757AC_0 vss vdd csvco_branch_2/vbp vdd csvco_branch_2/vbp
+ sky130_fd_pr__pfet_01v8_4757AC
Xcsvco_branch_0 vctrl out_vco csvco_branch_2/vbp D0 csvco_branch_1/in vss vdd csvco_branch
Xcsvco_branch_2 vctrl csvco_branch_2/in csvco_branch_2/vbp D0 out_vco vss vdd csvco_branch
Xcsvco_branch_1 vctrl csvco_branch_1/in csvco_branch_2/vbp D0 csvco_branch_2/in vss
+ vdd csvco_branch
.ends

.subckt ring_osc_buffer vss in_vco vdd o1 out_div out_pad
Xinverter_min_x4_1 vdd out_div vss out_pad inverter_min_x4
Xinverter_min_x4_0 vdd o1 vss out_div inverter_min_x4
Xinverter_min_x2_0 in_vco o1 vss vdd inverter_min_x2
.ends

.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X
X0 X B a_455_87# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 X a_194_125# a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_194_125# B a_158_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_158_392# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_355_368# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_194_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 a_455_87# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND B a_194_125# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X9 VGND a_194_125# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X
X0 VGND B a_143_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 X a_56_136# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VPWR B a_56_136# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_143_136# A a_56_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_56_136# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 X a_56_136# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__or2_1 A B VGND VNB VPB VPWR X
X0 VPWR A a_152_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_152_368# B a_63_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 X a_63_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 X a_63_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_63_368# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X5 VGND A a_63_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
.ends

.subckt div_by_5 nCLK vss vdd Q0 CLK nQ0 CLK_5 nQ2 Q1 Q1_shift
Xsky130_fd_sc_hs__xor2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_2/D sky130_fd_sc_hs__xor2_1
XDFlipFlop_0 vss nQ2 DFlipFlop_0/Q DFlipFlop_0/D vdd CLK nCLK DFlipFlop
XDFlipFlop_2 vss DFlipFlop_2/nQ Q1 DFlipFlop_2/D vdd CLK nCLK DFlipFlop
XDFlipFlop_1 vss nQ0 Q0 DFlipFlop_1/D vdd CLK nCLK DFlipFlop
XDFlipFlop_3 vss DFlipFlop_3/nQ Q1_shift Q1 vdd nCLK CLK DFlipFlop
Xsky130_fd_sc_hs__and2_1_0 Q1 Q0 vss vss vdd vdd DFlipFlop_0/D sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__and2_1_1 nQ2 nQ0 vss vss vdd vdd DFlipFlop_1/D sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__or2_1_0 Q1 Q1_shift vss vss vdd vdd CLK_5 sky130_fd_sc_hs__or2_1
.ends

.subckt sky130_fd_pr__nfet_01v8_AZESM8 a_n63_n151# a_n33_n125# a_n255_n151# a_33_n151#
+ a_n225_n125# a_63_n125# a_n129_n125# a_n159_n151# w_n455_n335# a_225_n151# a_255_n125#
+ a_129_n151# a_159_n125# a_n317_n125#
X0 a_159_n125# a_129_n151# a_63_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n225_n125# a_n255_n151# a_n317_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_63_n125# a_33_n151# a_n33_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_n129_n125# a_n159_n151# a_n225_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n33_n125# a_n63_n151# a_n129_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_255_n125# a_225_n151# a_159_n125# w_n455_n335# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_XJXT7S VSUBS a_n33_n125# a_n255_n154# a_33_n154# a_n225_n125#
+ a_n159_n154# a_63_n125# a_n129_n125# a_225_n154# a_129_n154# a_255_n125# a_159_n125#
+ a_n317_n125# w_n455_n344# a_n63_n154#
X0 a_n129_n125# a_n159_n154# a_n225_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X1 a_n33_n125# a_n63_n154# a_n129_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X2 a_255_n125# a_225_n154# a_159_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X3 a_159_n125# a_129_n154# a_63_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X4 a_n225_n125# a_n255_n154# a_n317_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
X5 a_63_n125# a_33_n154# a_n33_n125# w_n455_n344# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=150000u
.ends

.subckt inverter_cp_x2 in out vss vdd
Xsky130_fd_pr__nfet_01v8_AZESM8_0 in vss in in vss out out in vss in out in vss out
+ sky130_fd_pr__nfet_01v8_AZESM8
Xsky130_fd_pr__pfet_01v8_XJXT7S_0 vss vdd in in vdd in out out in in out vdd out vdd
+ in sky130_fd_pr__pfet_01v8_XJXT7S
.ends

.subckt pfd_cp_interface vss vdd Down QA QB nDown Up nUp
Xinverter_cp_x2_0 nDown Down vss vdd inverter_cp_x2
Xinverter_cp_x2_1 Up nUp vss vdd inverter_cp_x2
Xtrans_gate_0 nDown inverter_cp_x1_0/out vss vdd trans_gate
Xinverter_cp_x1_0 QB vss inverter_cp_x1_0/out vdd inverter_cp_x1
Xinverter_cp_x1_1 QA vss inverter_cp_x1_2/in vdd inverter_cp_x1
Xinverter_cp_x1_2 inverter_cp_x1_2/in vss Up vdd inverter_cp_x1
.ends

.subckt sky130_fd_pr__pfet_01v8_4F35BC VSUBS w_n359_n309# a_n63_n116# a_n159_n207#
+ a_n33_n90# a_n221_n90# a_159_n90#
X0 a_159_n90# a_n63_n116# a_63_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n129_n90# a_n159_n207# a_n221_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X2 a_63_n90# a_n159_n207# a_n33_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3 a_n33_n90# a_n63_n116# a_n129_n90# w_n359_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_C3YG4M a_n33_n45# a_33_n71# a_n129_71# w_n263_n255#
+ a_n125_n45# a_63_n45#
X0 a_63_n45# a_33_n71# a_n33_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n129_71# a_n125_n45# w_n263_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
.ends

.subckt nor_pfd out vss vdd A B
Xsky130_fd_pr__pfet_01v8_4F35BC_0 vss vdd B A out vdd vdd sky130_fd_pr__pfet_01v8_4F35BC
Xsky130_fd_pr__nfet_01v8_C3YG4M_0 out B A vss vss vss sky130_fd_pr__nfet_01v8_C3YG4M
.ends

.subckt dff_pfd vdd vss Q CLK Reset
Xnor_pfd_0 nor_pfd_2/A vss vdd CLK Q nor_pfd
Xnor_pfd_1 Q vss vdd nor_pfd_2/A nor_pfd_3/A nor_pfd
Xnor_pfd_2 nor_pfd_3/A vss vdd nor_pfd_2/A nor_pfd_2/B nor_pfd
Xnor_pfd_3 nor_pfd_2/B vss vdd nor_pfd_3/A Reset nor_pfd
.ends

.subckt sky130_fd_pr__nfet_01v8_ZCYAJJ w_n359_n255# a_n33_n45# a_n159_n173# a_n221_n45#
+ a_159_n45# a_n63_n71#
X0 a_63_n45# a_n159_n173# a_n33_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X1 a_n33_n45# a_n63_n71# a_n129_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X2 a_159_n45# a_n63_n71# a_63_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X3 a_n129_n45# a_n159_n173# a_n221_n45# w_n359_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_7T83YG VSUBS a_n125_n90# a_63_n90# a_33_n187# a_n99_n187#
+ a_n33_n90# w_n263_n309#
X0 a_63_n90# a_33_n187# a_n33_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X1 a_n33_n90# a_n99_n187# a_n125_n90# w_n263_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ZXAV3F a_n73_n45# a_n33_67# a_15_n45# w_n211_n255#
X0 a_15_n45# a_n33_67# a_n73_n45# w_n211_n255# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4F7GBC VSUBS a_n51_n187# a_n73_n90# a_15_n90# w_n211_n309#
X0 a_15_n90# a_n51_n187# a_n73_n90# w_n211_n309# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
.ends

.subckt and_pfd vss out vdd A B
Xsky130_fd_pr__nfet_01v8_ZCYAJJ_0 vss a_656_410# A vss vss B sky130_fd_pr__nfet_01v8_ZCYAJJ
Xsky130_fd_pr__pfet_01v8_7T83YG_0 vss vdd vdd B A a_656_410# vdd sky130_fd_pr__pfet_01v8_7T83YG
Xsky130_fd_pr__nfet_01v8_ZXAV3F_0 vss a_656_410# out vss sky130_fd_pr__nfet_01v8_ZXAV3F
Xsky130_fd_pr__pfet_01v8_4F7GBC_0 vss a_656_410# vdd out vdd sky130_fd_pr__pfet_01v8_4F7GBC
.ends

.subckt PFD vss vdd Down Up A B Reset
Xdff_pfd_0 vdd vss Up A Reset dff_pfd
Xdff_pfd_1 vdd vss Down B Reset dff_pfd
Xand_pfd_0 vss Reset vdd Up Down and_pfd
.ends

.subckt top_pll_v1 vdd in_ref w_13905_n238# vss vco_D0 iref_cp out_to_pad
Xloop_filter_0 lf_vc vco_vctrl vss loop_filter
Xcharge_pump_0 Down vco_vctrl iref_cp pswitch nDown biasp Up nswitch vss vdd nUp charge_pump
Xdiv_by_2_0 vss vdd out_by_2 n_out_by_2 out_buffer_div_2 out_to_div out_div_2 n_out_buffer_div_2
+ n_out_div_2 div_by_2
Xbuffer_salida_0 out_to_buffer out_to_pad vss vdd buffer_salida
Xring_osc_0 vco_vctrl vdd vss vco_D0 vco_out ring_osc
Xring_osc_buffer_0 vss vco_out vdd out_first_buffer out_to_div out_to_buffer ring_osc_buffer
Xdiv_by_5_0 n_out_by_2 vss vdd div_5_Q0 out_by_2 div_5_nQ0 out_div_by_5 div_5_nQ2
+ div_5_Q1 div_5_Q1_shift div_by_5
Xpfd_cp_interface_0 vss vdd Down QA QB nDown Up nUp pfd_cp_interface
XPFD_0 vss vdd QB QA in_ref out_div_by_5 pfd_reset PFD
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_2Y8F6P VSUBS c2_n3251_n3000# m4_n3351_n3100#
X0 c2_n3251_n3000# m4_n3351_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_8P223X VSUBS a_n2017_n1317# a_n1731_n1219# a_n1879_n1219#
+ a_n2017_n61# w_n2018_n202#
X0 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X1 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X2 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X3 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X4 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X5 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X6 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X7 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X8 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X9 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X10 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X11 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X12 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X13 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X14 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X15 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X16 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X17 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X18 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X19 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X20 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X21 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X22 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X23 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X24 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X25 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X26 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X27 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X28 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X29 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X30 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X31 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X32 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X33 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X34 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X35 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X36 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X37 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X38 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X39 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X40 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X41 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X42 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X43 a_n1879_n1219# a_n2017_n1317# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X44 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X45 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X46 a_n1731_n1219# a_n2017_n61# w_n2018_n202# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X47 w_n2018_n202# a_n2017_n61# a_n1731_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X48 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
X49 a_n1731_n1219# a_n2017_n1317# a_n1879_n1219# w_n2018_n202# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=450000u
.ends

.subckt bias VSUBS vdd iref_0 iref_1 iref_2 iref_5 iref_6 iref_7 iref_8 iref_9 iref
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_5 VSUBS iref m1_20168_984# iref m1_20168_984#
+ vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_6 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_6/a_n1731_n1219#
+ iref_5 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_7 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_7/a_n1731_n1219#
+ iref_6 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_9 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_9/a_n1731_n1219#
+ iref_8 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_8 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_8/a_n1731_n1219#
+ iref_7 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_10 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_10/a_n1731_n1219#
+ iref_9 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_0 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_0/a_n1731_n1219#
+ iref_0 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_1 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_1/a_n1731_n1219#
+ iref_1 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_2 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_2/a_n1731_n1219#
+ iref_2 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_3 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_3/a_n1731_n1219#
+ iref_3 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
Xsky130_fd_pr__pfet_01v8_lvt_8P223X_4 VSUBS iref sky130_fd_pr__pfet_01v8_lvt_8P223X_4/a_n1731_n1219#
+ iref_4 m1_20168_984# vdd sky130_fd_pr__pfet_01v8_lvt_8P223X
.ends

.subckt mimcap_decoup_1x5 VSUBS t b
Xdecap[0] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[1] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[2] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[3] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xdecap[4] VSUBS t b sky130_fd_pr__cap_mim_m3_2_2Y8F6P
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WHJTNJ VSUBS m3_n4309_50# m3_n4309_n4250# c1_n4209_n4150#
+ c1_110_n4150# m3_10_n4250#
X0 c1_n4209_n4150# m3_n4309_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X1 c1_110_n4150# m3_10_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X2 c1_n4209_n4150# m3_n4309_50# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
X3 c1_110_n4150# m3_10_n4250# sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2e+07u
.ends

.subckt cap3_loop_filter VSUBS in out
Xsky130_fd_pr__cap_mim_m3_1_WHJTNJ_0 VSUBS out out in in out sky130_fd_pr__cap_mim_m3_1_WHJTNJ
.ends

.subckt sky130_fd_pr__nfet_01v8_U2JGXT w_n226_n510# a_n118_n388# a_n88_n300# a_30_n300#
X0 a_30_n300# a_n118_n388# a_n88_n300# w_n226_n510# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
.ends

.subckt loop_filter_v2 vc_pex D0_cap in vss
Xcap1_loop_filter_0 vss vc_pex vss cap1_loop_filter
Xcap3_loop_filter_0 vss cap3_loop_filter_0/in vss cap3_loop_filter
Xcap2_loop_filter_0 vss in vss cap2_loop_filter
Xsky130_fd_pr__nfet_01v8_U2JGXT_0 vss D0_cap in cap3_loop_filter_0/in sky130_fd_pr__nfet_01v8_U2JGXT
Xres_loop_filter_0 vss res_loop_filter_2/out in res_loop_filter
Xres_loop_filter_1 vss res_loop_filter_2/out vc_pex res_loop_filter
Xres_loop_filter_2 vss res_loop_filter_2/out vc_pex res_loop_filter
.ends

.subckt top_pll_v2 vdd in_ref w_13905_n238# vss D0_vco iref_cp DO_cap out_to_pad
Xcharge_pump_0 Down vco_vctrl iref_cp pswitch nDown biasp Up nswitch vss vdd nUp charge_pump
Xloop_filter_v2_0 lf_vc DO_cap vco_vctrl vss loop_filter_v2
Xdiv_by_2_0 vss vdd out_by_2 n_out_by_2 out_buffer_div_2 out_to_div out_div_2 n_out_buffer_div_2
+ n_out_div_2 div_by_2
Xbuffer_salida_0 out_to_buffer out_to_pad vss vdd buffer_salida
Xring_osc_0 vco_vctrl vdd vss D0_vco vco_out ring_osc
Xring_osc_buffer_0 vss vco_out vdd out_first_buffer out_to_div out_to_buffer ring_osc_buffer
Xdiv_by_5_0 n_out_by_2 vss vdd div_5_Q0 out_by_2 div_5_nQ0 out_div_by_5 div_5_nQ2
+ div_5_Q1 div_5_Q1_shift div_by_5
Xpfd_cp_interface_0 vss vdd Down QA QB nDown Up nUp pfd_cp_interface
XPFD_0 vss vdd QB QA in_ref out_div_by_5 pfd_reset PFD
.ends

*.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
*+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
*+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
*+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
*+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
*+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
*+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
*+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
*+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[2] io_clamp_low[0] io_clamp_low[2]
*+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
*+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
*+ io_in[26] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9]
*+ io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12] io_in_3v3[13] io_in_3v3[14]
*+ io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18] io_in_3v3[19] io_in_3v3[1]
*+ io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23] io_in_3v3[24] io_in_3v3[25]
*+ io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4] io_in_3v3[5] io_in_3v3[6] io_in_3v3[7]
*+ io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
*+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
*+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[2] io_oeb[3]
*+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
*+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
*+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
*+ io_out[26] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8]
*+ io_out[9] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
*+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
*+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
*+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
*+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
*+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
*+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
*+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
*+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
*+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
*+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
*+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
*+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
*+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
*+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
*+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
*+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
*+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
*+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
*+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
*+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
*+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
*+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
*+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
*+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
*+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
*+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
*+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
*+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
*+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
*+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
*+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
*+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
*+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
*+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
*+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
*+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
*+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
*+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
*+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
*+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
*+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
*+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
*+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
*+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
*+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
*+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
*+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
*+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
*+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
*+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
*+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
*+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
*+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
*+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
*+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
*+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
*+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
*+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
*+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
*+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
*+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
*+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
*+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
*+ user_clock2 user_irq[0] user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2
*+ vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
*+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
*+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
*+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
*+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
*+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
*+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
*+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
*+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
*+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
*+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
*+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
*+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
*+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
*+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
*+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
*+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xres_amp_top_0 bias_0/iref_9 bias_0/iref_8 vssa1 bias_0/iref_6 bias_0/iref_7 bias_0/iref_5
+ vdda1 io_analog[6] gpio_noesd[4] gpio_noesd[5] gpio_noesd[6] gpio_noesd[3] gpio_noesd[2]
+ io_analog[2] io_analog[0] gpio_noesd[1] io_analog[1] io_analog[3] io_analog[4] res_amp_top
Xtop_pll_v1_0 vdda1 io_analog[10] vssa1 vssa1 gpio_noesd[7] bias_0/iref_2 io_analog[9]
+ top_pll_v1
Xtop_pll_v1_1 vdda1 io_analog[10] vssa1 vssa1 gpio_noesd[7] bias_0/iref_0 io_analog[7]
+ top_pll_v1
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[0] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[1] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[2] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[3] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[4] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[5] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[6] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[7] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_0[8] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xbias_0 vssa1 vdda1 bias_0/iref_0 bias_0/iref_1 bias_0/iref_2 bias_0/iref_5 bias_0/iref_6
+ bias_0/iref_7 bias_0/iref_8 bias_0/iref_9 io_analog[5] bias
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[0] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[1] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[2] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[3] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[4] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[5] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[6] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[7] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_1[8] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xmimcap_decoup_1x5_0[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_0[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_0[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_1[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_1[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_1[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[0] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[1] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[2] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[3] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[4] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[5] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xsky130_fd_pr__cap_mim_m3_2_2Y8F6P_2[6] vssa1 vdda1 vssa1 sky130_fd_pr__cap_mim_m3_2_2Y8F6P
Xmimcap_decoup_1x5_2[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_2[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_2[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_3[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_3[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_3[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_4[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_4[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_4[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_5[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_5[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_5[2] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_6[0] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xmimcap_decoup_1x5_6[1] vssa1 vdda1 vssa1 mimcap_decoup_1x5
Xtop_pll_v2_0 vdda1 io_analog[10] vssa1 vssa1 gpio_noesd[7] bias_0/iref_1 gpio_noesd[8]
+ io_analog[8] top_pll_v2
.end

