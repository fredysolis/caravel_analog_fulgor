magic
tech sky130A
magscale 1 2
timestamp 1623991863
<< error_p >>
rect -1887 331 -1857 335
rect -1791 331 -1761 335
rect -1695 331 -1665 335
rect -1599 331 -1569 335
rect -1503 331 -1473 335
rect -1407 331 -1377 335
rect -1311 331 -1281 335
rect -1215 331 -1185 335
rect -1119 331 -1089 335
rect -1023 331 -993 335
rect -927 331 -897 335
rect -831 331 -801 335
rect -735 331 -705 335
rect -639 331 -609 335
rect -543 331 -513 335
rect -447 331 -417 335
rect -351 331 -321 335
rect -255 331 -225 335
rect -159 331 -129 335
rect -63 331 -33 335
rect 33 331 63 335
rect 129 331 159 335
rect 225 331 255 335
rect 321 331 351 335
rect 417 331 447 335
rect 513 331 543 335
rect 609 331 639 335
rect 705 331 735 335
rect 801 331 831 335
rect 897 331 927 335
rect 993 331 1023 335
rect 1089 331 1119 335
rect 1185 331 1215 335
rect 1281 331 1311 335
rect 1377 331 1407 335
rect 1473 331 1503 335
rect 1569 331 1599 335
rect 1665 331 1695 335
rect 1761 331 1791 335
rect -1887 -335 -1857 -331
rect -1791 -335 -1761 -331
rect -1695 -335 -1665 -331
rect -1599 -335 -1569 -331
rect -1503 -335 -1473 -331
rect -1407 -335 -1377 -331
rect -1311 -335 -1281 -331
rect -1215 -335 -1185 -331
rect -1119 -335 -1089 -331
rect -1023 -335 -993 -331
rect -927 -335 -897 -331
rect -831 -335 -801 -331
rect -735 -335 -705 -331
rect -639 -335 -609 -331
rect -543 -335 -513 -331
rect -447 -335 -417 -331
rect -351 -335 -321 -331
rect -255 -335 -225 -331
rect -159 -335 -129 -331
rect -63 -335 -33 -331
rect 33 -335 63 -331
rect 129 -335 159 -331
rect 225 -335 255 -331
rect 321 -335 351 -331
rect 417 -335 447 -331
rect 513 -335 543 -331
rect 609 -335 639 -331
rect 705 -335 735 -331
rect 801 -335 831 -331
rect 897 -335 927 -331
rect 993 -335 1023 -331
rect 1089 -335 1119 -331
rect 1185 -335 1215 -331
rect 1281 -335 1311 -331
rect 1377 -335 1407 -331
rect 1473 -335 1503 -331
rect 1569 -335 1599 -331
rect 1665 -335 1695 -331
rect 1761 -335 1791 -331
<< pwell >>
rect -2087 -519 2087 519
<< nmoslvt >>
rect -1887 109 -1857 309
rect -1791 109 -1761 309
rect -1695 109 -1665 309
rect -1599 109 -1569 309
rect -1503 109 -1473 309
rect -1407 109 -1377 309
rect -1311 109 -1281 309
rect -1215 109 -1185 309
rect -1119 109 -1089 309
rect -1023 109 -993 309
rect -927 109 -897 309
rect -831 109 -801 309
rect -735 109 -705 309
rect -639 109 -609 309
rect -543 109 -513 309
rect -447 109 -417 309
rect -351 109 -321 309
rect -255 109 -225 309
rect -159 109 -129 309
rect -63 109 -33 309
rect 33 109 63 309
rect 129 109 159 309
rect 225 109 255 309
rect 321 109 351 309
rect 417 109 447 309
rect 513 109 543 309
rect 609 109 639 309
rect 705 109 735 309
rect 801 109 831 309
rect 897 109 927 309
rect 993 109 1023 309
rect 1089 109 1119 309
rect 1185 109 1215 309
rect 1281 109 1311 309
rect 1377 109 1407 309
rect 1473 109 1503 309
rect 1569 109 1599 309
rect 1665 109 1695 309
rect 1761 109 1791 309
rect 1857 109 1887 309
rect -1887 -309 -1857 -109
rect -1791 -309 -1761 -109
rect -1695 -309 -1665 -109
rect -1599 -309 -1569 -109
rect -1503 -309 -1473 -109
rect -1407 -309 -1377 -109
rect -1311 -309 -1281 -109
rect -1215 -309 -1185 -109
rect -1119 -309 -1089 -109
rect -1023 -309 -993 -109
rect -927 -309 -897 -109
rect -831 -309 -801 -109
rect -735 -309 -705 -109
rect -639 -309 -609 -109
rect -543 -309 -513 -109
rect -447 -309 -417 -109
rect -351 -309 -321 -109
rect -255 -309 -225 -109
rect -159 -309 -129 -109
rect -63 -309 -33 -109
rect 33 -309 63 -109
rect 129 -309 159 -109
rect 225 -309 255 -109
rect 321 -309 351 -109
rect 417 -309 447 -109
rect 513 -309 543 -109
rect 609 -309 639 -109
rect 705 -309 735 -109
rect 801 -309 831 -109
rect 897 -309 927 -109
rect 993 -309 1023 -109
rect 1089 -309 1119 -109
rect 1185 -309 1215 -109
rect 1281 -309 1311 -109
rect 1377 -309 1407 -109
rect 1473 -309 1503 -109
rect 1569 -309 1599 -109
rect 1665 -309 1695 -109
rect 1761 -309 1791 -109
rect 1857 -309 1887 -109
<< ndiff >>
rect -1949 297 -1887 309
rect -1949 121 -1937 297
rect -1903 121 -1887 297
rect -1949 109 -1887 121
rect -1857 297 -1791 309
rect -1857 121 -1841 297
rect -1807 121 -1791 297
rect -1857 109 -1791 121
rect -1761 297 -1695 309
rect -1761 121 -1745 297
rect -1711 121 -1695 297
rect -1761 109 -1695 121
rect -1665 297 -1599 309
rect -1665 121 -1649 297
rect -1615 121 -1599 297
rect -1665 109 -1599 121
rect -1569 297 -1503 309
rect -1569 121 -1553 297
rect -1519 121 -1503 297
rect -1569 109 -1503 121
rect -1473 297 -1407 309
rect -1473 121 -1457 297
rect -1423 121 -1407 297
rect -1473 109 -1407 121
rect -1377 297 -1311 309
rect -1377 121 -1361 297
rect -1327 121 -1311 297
rect -1377 109 -1311 121
rect -1281 297 -1215 309
rect -1281 121 -1265 297
rect -1231 121 -1215 297
rect -1281 109 -1215 121
rect -1185 297 -1119 309
rect -1185 121 -1169 297
rect -1135 121 -1119 297
rect -1185 109 -1119 121
rect -1089 297 -1023 309
rect -1089 121 -1073 297
rect -1039 121 -1023 297
rect -1089 109 -1023 121
rect -993 297 -927 309
rect -993 121 -977 297
rect -943 121 -927 297
rect -993 109 -927 121
rect -897 297 -831 309
rect -897 121 -881 297
rect -847 121 -831 297
rect -897 109 -831 121
rect -801 297 -735 309
rect -801 121 -785 297
rect -751 121 -735 297
rect -801 109 -735 121
rect -705 297 -639 309
rect -705 121 -689 297
rect -655 121 -639 297
rect -705 109 -639 121
rect -609 297 -543 309
rect -609 121 -593 297
rect -559 121 -543 297
rect -609 109 -543 121
rect -513 297 -447 309
rect -513 121 -497 297
rect -463 121 -447 297
rect -513 109 -447 121
rect -417 297 -351 309
rect -417 121 -401 297
rect -367 121 -351 297
rect -417 109 -351 121
rect -321 297 -255 309
rect -321 121 -305 297
rect -271 121 -255 297
rect -321 109 -255 121
rect -225 297 -159 309
rect -225 121 -209 297
rect -175 121 -159 297
rect -225 109 -159 121
rect -129 297 -63 309
rect -129 121 -113 297
rect -79 121 -63 297
rect -129 109 -63 121
rect -33 297 33 309
rect -33 121 -17 297
rect 17 121 33 297
rect -33 109 33 121
rect 63 297 129 309
rect 63 121 79 297
rect 113 121 129 297
rect 63 109 129 121
rect 159 297 225 309
rect 159 121 175 297
rect 209 121 225 297
rect 159 109 225 121
rect 255 297 321 309
rect 255 121 271 297
rect 305 121 321 297
rect 255 109 321 121
rect 351 297 417 309
rect 351 121 367 297
rect 401 121 417 297
rect 351 109 417 121
rect 447 297 513 309
rect 447 121 463 297
rect 497 121 513 297
rect 447 109 513 121
rect 543 297 609 309
rect 543 121 559 297
rect 593 121 609 297
rect 543 109 609 121
rect 639 297 705 309
rect 639 121 655 297
rect 689 121 705 297
rect 639 109 705 121
rect 735 297 801 309
rect 735 121 751 297
rect 785 121 801 297
rect 735 109 801 121
rect 831 297 897 309
rect 831 121 847 297
rect 881 121 897 297
rect 831 109 897 121
rect 927 297 993 309
rect 927 121 943 297
rect 977 121 993 297
rect 927 109 993 121
rect 1023 297 1089 309
rect 1023 121 1039 297
rect 1073 121 1089 297
rect 1023 109 1089 121
rect 1119 297 1185 309
rect 1119 121 1135 297
rect 1169 121 1185 297
rect 1119 109 1185 121
rect 1215 297 1281 309
rect 1215 121 1231 297
rect 1265 121 1281 297
rect 1215 109 1281 121
rect 1311 297 1377 309
rect 1311 121 1327 297
rect 1361 121 1377 297
rect 1311 109 1377 121
rect 1407 297 1473 309
rect 1407 121 1423 297
rect 1457 121 1473 297
rect 1407 109 1473 121
rect 1503 297 1569 309
rect 1503 121 1519 297
rect 1553 121 1569 297
rect 1503 109 1569 121
rect 1599 297 1665 309
rect 1599 121 1615 297
rect 1649 121 1665 297
rect 1599 109 1665 121
rect 1695 297 1761 309
rect 1695 121 1711 297
rect 1745 121 1761 297
rect 1695 109 1761 121
rect 1791 297 1857 309
rect 1791 121 1807 297
rect 1841 121 1857 297
rect 1791 109 1857 121
rect 1887 297 1949 309
rect 1887 121 1903 297
rect 1937 121 1949 297
rect 1887 109 1949 121
rect -1949 -121 -1887 -109
rect -1949 -297 -1937 -121
rect -1903 -297 -1887 -121
rect -1949 -309 -1887 -297
rect -1857 -121 -1791 -109
rect -1857 -297 -1841 -121
rect -1807 -297 -1791 -121
rect -1857 -309 -1791 -297
rect -1761 -121 -1695 -109
rect -1761 -297 -1745 -121
rect -1711 -297 -1695 -121
rect -1761 -309 -1695 -297
rect -1665 -121 -1599 -109
rect -1665 -297 -1649 -121
rect -1615 -297 -1599 -121
rect -1665 -309 -1599 -297
rect -1569 -121 -1503 -109
rect -1569 -297 -1553 -121
rect -1519 -297 -1503 -121
rect -1569 -309 -1503 -297
rect -1473 -121 -1407 -109
rect -1473 -297 -1457 -121
rect -1423 -297 -1407 -121
rect -1473 -309 -1407 -297
rect -1377 -121 -1311 -109
rect -1377 -297 -1361 -121
rect -1327 -297 -1311 -121
rect -1377 -309 -1311 -297
rect -1281 -121 -1215 -109
rect -1281 -297 -1265 -121
rect -1231 -297 -1215 -121
rect -1281 -309 -1215 -297
rect -1185 -121 -1119 -109
rect -1185 -297 -1169 -121
rect -1135 -297 -1119 -121
rect -1185 -309 -1119 -297
rect -1089 -121 -1023 -109
rect -1089 -297 -1073 -121
rect -1039 -297 -1023 -121
rect -1089 -309 -1023 -297
rect -993 -121 -927 -109
rect -993 -297 -977 -121
rect -943 -297 -927 -121
rect -993 -309 -927 -297
rect -897 -121 -831 -109
rect -897 -297 -881 -121
rect -847 -297 -831 -121
rect -897 -309 -831 -297
rect -801 -121 -735 -109
rect -801 -297 -785 -121
rect -751 -297 -735 -121
rect -801 -309 -735 -297
rect -705 -121 -639 -109
rect -705 -297 -689 -121
rect -655 -297 -639 -121
rect -705 -309 -639 -297
rect -609 -121 -543 -109
rect -609 -297 -593 -121
rect -559 -297 -543 -121
rect -609 -309 -543 -297
rect -513 -121 -447 -109
rect -513 -297 -497 -121
rect -463 -297 -447 -121
rect -513 -309 -447 -297
rect -417 -121 -351 -109
rect -417 -297 -401 -121
rect -367 -297 -351 -121
rect -417 -309 -351 -297
rect -321 -121 -255 -109
rect -321 -297 -305 -121
rect -271 -297 -255 -121
rect -321 -309 -255 -297
rect -225 -121 -159 -109
rect -225 -297 -209 -121
rect -175 -297 -159 -121
rect -225 -309 -159 -297
rect -129 -121 -63 -109
rect -129 -297 -113 -121
rect -79 -297 -63 -121
rect -129 -309 -63 -297
rect -33 -121 33 -109
rect -33 -297 -17 -121
rect 17 -297 33 -121
rect -33 -309 33 -297
rect 63 -121 129 -109
rect 63 -297 79 -121
rect 113 -297 129 -121
rect 63 -309 129 -297
rect 159 -121 225 -109
rect 159 -297 175 -121
rect 209 -297 225 -121
rect 159 -309 225 -297
rect 255 -121 321 -109
rect 255 -297 271 -121
rect 305 -297 321 -121
rect 255 -309 321 -297
rect 351 -121 417 -109
rect 351 -297 367 -121
rect 401 -297 417 -121
rect 351 -309 417 -297
rect 447 -121 513 -109
rect 447 -297 463 -121
rect 497 -297 513 -121
rect 447 -309 513 -297
rect 543 -121 609 -109
rect 543 -297 559 -121
rect 593 -297 609 -121
rect 543 -309 609 -297
rect 639 -121 705 -109
rect 639 -297 655 -121
rect 689 -297 705 -121
rect 639 -309 705 -297
rect 735 -121 801 -109
rect 735 -297 751 -121
rect 785 -297 801 -121
rect 735 -309 801 -297
rect 831 -121 897 -109
rect 831 -297 847 -121
rect 881 -297 897 -121
rect 831 -309 897 -297
rect 927 -121 993 -109
rect 927 -297 943 -121
rect 977 -297 993 -121
rect 927 -309 993 -297
rect 1023 -121 1089 -109
rect 1023 -297 1039 -121
rect 1073 -297 1089 -121
rect 1023 -309 1089 -297
rect 1119 -121 1185 -109
rect 1119 -297 1135 -121
rect 1169 -297 1185 -121
rect 1119 -309 1185 -297
rect 1215 -121 1281 -109
rect 1215 -297 1231 -121
rect 1265 -297 1281 -121
rect 1215 -309 1281 -297
rect 1311 -121 1377 -109
rect 1311 -297 1327 -121
rect 1361 -297 1377 -121
rect 1311 -309 1377 -297
rect 1407 -121 1473 -109
rect 1407 -297 1423 -121
rect 1457 -297 1473 -121
rect 1407 -309 1473 -297
rect 1503 -121 1569 -109
rect 1503 -297 1519 -121
rect 1553 -297 1569 -121
rect 1503 -309 1569 -297
rect 1599 -121 1665 -109
rect 1599 -297 1615 -121
rect 1649 -297 1665 -121
rect 1599 -309 1665 -297
rect 1695 -121 1761 -109
rect 1695 -297 1711 -121
rect 1745 -297 1761 -121
rect 1695 -309 1761 -297
rect 1791 -121 1857 -109
rect 1791 -297 1807 -121
rect 1841 -297 1857 -121
rect 1791 -309 1857 -297
rect 1887 -121 1949 -109
rect 1887 -297 1903 -121
rect 1937 -297 1949 -121
rect 1887 -309 1949 -297
<< ndiffc >>
rect -1937 121 -1903 297
rect -1841 121 -1807 297
rect -1745 121 -1711 297
rect -1649 121 -1615 297
rect -1553 121 -1519 297
rect -1457 121 -1423 297
rect -1361 121 -1327 297
rect -1265 121 -1231 297
rect -1169 121 -1135 297
rect -1073 121 -1039 297
rect -977 121 -943 297
rect -881 121 -847 297
rect -785 121 -751 297
rect -689 121 -655 297
rect -593 121 -559 297
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect 559 121 593 297
rect 655 121 689 297
rect 751 121 785 297
rect 847 121 881 297
rect 943 121 977 297
rect 1039 121 1073 297
rect 1135 121 1169 297
rect 1231 121 1265 297
rect 1327 121 1361 297
rect 1423 121 1457 297
rect 1519 121 1553 297
rect 1615 121 1649 297
rect 1711 121 1745 297
rect 1807 121 1841 297
rect 1903 121 1937 297
rect -1937 -297 -1903 -121
rect -1841 -297 -1807 -121
rect -1745 -297 -1711 -121
rect -1649 -297 -1615 -121
rect -1553 -297 -1519 -121
rect -1457 -297 -1423 -121
rect -1361 -297 -1327 -121
rect -1265 -297 -1231 -121
rect -1169 -297 -1135 -121
rect -1073 -297 -1039 -121
rect -977 -297 -943 -121
rect -881 -297 -847 -121
rect -785 -297 -751 -121
rect -689 -297 -655 -121
rect -593 -297 -559 -121
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect 559 -297 593 -121
rect 655 -297 689 -121
rect 751 -297 785 -121
rect 847 -297 881 -121
rect 943 -297 977 -121
rect 1039 -297 1073 -121
rect 1135 -297 1169 -121
rect 1231 -297 1265 -121
rect 1327 -297 1361 -121
rect 1423 -297 1457 -121
rect 1519 -297 1553 -121
rect 1615 -297 1649 -121
rect 1711 -297 1745 -121
rect 1807 -297 1841 -121
rect 1903 -297 1937 -121
<< psubdiff >>
rect -2051 449 -1955 483
rect 1955 449 2051 483
rect 2017 387 2051 449
rect 2017 -449 2051 -387
rect -2051 -483 -1955 -449
rect 1955 -483 2051 -449
<< psubdiffcont >>
rect -1955 449 1955 483
rect 2017 -387 2051 387
rect -1955 -483 1955 -449
<< poly >>
rect -1887 309 -1857 331
rect -1791 309 -1761 331
rect -1695 309 -1665 331
rect -1599 309 -1569 331
rect -1503 309 -1473 331
rect -1407 309 -1377 331
rect -1311 309 -1281 331
rect -1215 309 -1185 331
rect -1119 309 -1089 331
rect -1023 309 -993 331
rect -927 309 -897 331
rect -831 309 -801 331
rect -735 309 -705 331
rect -639 309 -609 331
rect -543 309 -513 331
rect -447 309 -417 331
rect -351 309 -321 331
rect -255 309 -225 331
rect -159 309 -129 331
rect -63 309 -33 331
rect 33 309 63 331
rect 129 309 159 331
rect 225 309 255 331
rect 321 309 351 331
rect 417 309 447 331
rect 513 309 543 331
rect 609 309 639 331
rect 705 309 735 331
rect 801 309 831 331
rect 897 309 927 331
rect 993 309 1023 331
rect 1089 309 1119 331
rect 1185 309 1215 331
rect 1281 309 1311 331
rect 1377 309 1407 331
rect 1473 309 1503 331
rect 1569 309 1599 331
rect 1665 309 1695 331
rect 1761 309 1791 331
rect 1857 309 1887 335
rect -1887 87 -1857 109
rect -1791 87 -1761 109
rect -1695 87 -1665 109
rect -1599 87 -1569 109
rect -1503 87 -1473 109
rect -1407 87 -1377 109
rect -1311 87 -1281 109
rect -1215 87 -1185 109
rect -1119 87 -1089 109
rect -1023 87 -993 109
rect -927 87 -897 109
rect -831 87 -801 109
rect -735 87 -705 109
rect -639 87 -609 109
rect -543 87 -513 109
rect -447 87 -417 109
rect -351 87 -321 109
rect -255 87 -225 109
rect -159 87 -129 109
rect -63 87 -33 109
rect 33 87 63 109
rect 129 87 159 109
rect 225 87 255 109
rect 321 87 351 109
rect 417 87 447 109
rect 513 87 543 109
rect 609 87 639 109
rect 705 87 735 109
rect 801 87 831 109
rect 897 87 927 109
rect 993 87 1023 109
rect 1089 87 1119 109
rect 1185 87 1215 109
rect 1281 87 1311 109
rect 1377 87 1407 109
rect 1473 87 1503 109
rect 1569 87 1599 109
rect 1665 87 1695 109
rect 1761 87 1791 109
rect 1857 87 1887 109
rect -1905 -87 1905 87
rect -1887 -109 -1857 -87
rect -1791 -109 -1761 -87
rect -1695 -109 -1665 -87
rect -1599 -109 -1569 -87
rect -1503 -109 -1473 -87
rect -1407 -109 -1377 -87
rect -1311 -109 -1281 -87
rect -1215 -109 -1185 -87
rect -1119 -109 -1089 -87
rect -1023 -109 -993 -87
rect -927 -109 -897 -87
rect -831 -109 -801 -87
rect -735 -109 -705 -87
rect -639 -109 -609 -87
rect -543 -109 -513 -87
rect -447 -109 -417 -87
rect -351 -109 -321 -87
rect -255 -109 -225 -87
rect -159 -109 -129 -87
rect -63 -109 -33 -87
rect 33 -109 63 -87
rect 129 -109 159 -87
rect 225 -109 255 -87
rect 321 -109 351 -87
rect 417 -109 447 -87
rect 513 -109 543 -87
rect 609 -109 639 -87
rect 705 -109 735 -87
rect 801 -109 831 -87
rect 897 -109 927 -87
rect 993 -109 1023 -87
rect 1089 -109 1119 -87
rect 1185 -109 1215 -87
rect 1281 -109 1311 -87
rect 1377 -109 1407 -87
rect 1473 -109 1503 -87
rect 1569 -109 1599 -87
rect 1665 -109 1695 -87
rect 1761 -109 1791 -87
rect 1857 -109 1887 -87
rect -1887 -331 -1857 -309
rect -1791 -331 -1761 -309
rect -1695 -331 -1665 -309
rect -1599 -331 -1569 -309
rect -1503 -331 -1473 -309
rect -1407 -331 -1377 -309
rect -1311 -331 -1281 -309
rect -1215 -331 -1185 -309
rect -1119 -331 -1089 -309
rect -1023 -331 -993 -309
rect -927 -331 -897 -309
rect -831 -331 -801 -309
rect -735 -331 -705 -309
rect -639 -331 -609 -309
rect -543 -331 -513 -309
rect -447 -331 -417 -309
rect -351 -331 -321 -309
rect -255 -331 -225 -309
rect -159 -331 -129 -309
rect -63 -331 -33 -309
rect 33 -331 63 -309
rect 129 -331 159 -309
rect 225 -331 255 -309
rect 321 -331 351 -309
rect 417 -331 447 -309
rect 513 -331 543 -309
rect 609 -331 639 -309
rect 705 -331 735 -309
rect 801 -331 831 -309
rect 897 -331 927 -309
rect 993 -331 1023 -309
rect 1089 -331 1119 -309
rect 1185 -331 1215 -309
rect 1281 -331 1311 -309
rect 1377 -331 1407 -309
rect 1473 -331 1503 -309
rect 1569 -331 1599 -309
rect 1665 -331 1695 -309
rect 1761 -331 1791 -309
rect 1857 -335 1887 -309
<< locali >>
rect -2051 449 -1955 483
rect 1955 449 2051 483
rect 2017 387 2051 449
rect -1937 297 -1903 313
rect -1937 105 -1903 121
rect -1841 297 -1807 313
rect -1841 105 -1807 121
rect -1745 297 -1711 313
rect -1745 105 -1711 121
rect -1649 297 -1615 313
rect -1649 105 -1615 121
rect -1553 297 -1519 313
rect -1553 105 -1519 121
rect -1457 297 -1423 313
rect -1457 105 -1423 121
rect -1361 297 -1327 313
rect -1361 105 -1327 121
rect -1265 297 -1231 313
rect -1265 105 -1231 121
rect -1169 297 -1135 313
rect -1169 105 -1135 121
rect -1073 297 -1039 313
rect -1073 105 -1039 121
rect -977 297 -943 313
rect -977 105 -943 121
rect -881 297 -847 313
rect -881 105 -847 121
rect -785 297 -751 313
rect -785 105 -751 121
rect -689 297 -655 313
rect -689 105 -655 121
rect -593 297 -559 313
rect -593 105 -559 121
rect -497 297 -463 313
rect -497 105 -463 121
rect -401 297 -367 313
rect -401 105 -367 121
rect -305 297 -271 313
rect -305 105 -271 121
rect -209 297 -175 313
rect -209 105 -175 121
rect -113 297 -79 313
rect -113 105 -79 121
rect -17 297 17 313
rect -17 105 17 121
rect 79 297 113 313
rect 79 105 113 121
rect 175 297 209 313
rect 175 105 209 121
rect 271 297 305 313
rect 271 105 305 121
rect 367 297 401 313
rect 367 105 401 121
rect 463 297 497 313
rect 463 105 497 121
rect 559 297 593 313
rect 559 105 593 121
rect 655 297 689 313
rect 655 105 689 121
rect 751 297 785 313
rect 751 105 785 121
rect 847 297 881 313
rect 847 105 881 121
rect 943 297 977 313
rect 943 105 977 121
rect 1039 297 1073 313
rect 1039 105 1073 121
rect 1135 297 1169 313
rect 1135 105 1169 121
rect 1231 297 1265 313
rect 1231 105 1265 121
rect 1327 297 1361 313
rect 1327 105 1361 121
rect 1423 297 1457 313
rect 1423 105 1457 121
rect 1519 297 1553 313
rect 1519 105 1553 121
rect 1615 297 1649 313
rect 1615 105 1649 121
rect 1711 297 1745 313
rect 1711 105 1745 121
rect 1807 297 1841 313
rect 1807 105 1841 121
rect 1903 297 1937 313
rect 1903 105 1937 121
rect -1937 -121 -1903 -105
rect -1937 -313 -1903 -297
rect -1841 -121 -1807 -105
rect -1841 -313 -1807 -297
rect -1745 -121 -1711 -105
rect -1745 -313 -1711 -297
rect -1649 -121 -1615 -105
rect -1649 -313 -1615 -297
rect -1553 -121 -1519 -105
rect -1553 -313 -1519 -297
rect -1457 -121 -1423 -105
rect -1457 -313 -1423 -297
rect -1361 -121 -1327 -105
rect -1361 -313 -1327 -297
rect -1265 -121 -1231 -105
rect -1265 -313 -1231 -297
rect -1169 -121 -1135 -105
rect -1169 -313 -1135 -297
rect -1073 -121 -1039 -105
rect -1073 -313 -1039 -297
rect -977 -121 -943 -105
rect -977 -313 -943 -297
rect -881 -121 -847 -105
rect -881 -313 -847 -297
rect -785 -121 -751 -105
rect -785 -313 -751 -297
rect -689 -121 -655 -105
rect -689 -313 -655 -297
rect -593 -121 -559 -105
rect -593 -313 -559 -297
rect -497 -121 -463 -105
rect -497 -313 -463 -297
rect -401 -121 -367 -105
rect -401 -313 -367 -297
rect -305 -121 -271 -105
rect -305 -313 -271 -297
rect -209 -121 -175 -105
rect -209 -313 -175 -297
rect -113 -121 -79 -105
rect -113 -313 -79 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 79 -121 113 -105
rect 79 -313 113 -297
rect 175 -121 209 -105
rect 175 -313 209 -297
rect 271 -121 305 -105
rect 271 -313 305 -297
rect 367 -121 401 -105
rect 367 -313 401 -297
rect 463 -121 497 -105
rect 463 -313 497 -297
rect 559 -121 593 -105
rect 559 -313 593 -297
rect 655 -121 689 -105
rect 655 -313 689 -297
rect 751 -121 785 -105
rect 751 -313 785 -297
rect 847 -121 881 -105
rect 847 -313 881 -297
rect 943 -121 977 -105
rect 943 -313 977 -297
rect 1039 -121 1073 -105
rect 1039 -313 1073 -297
rect 1135 -121 1169 -105
rect 1135 -313 1169 -297
rect 1231 -121 1265 -105
rect 1231 -313 1265 -297
rect 1327 -121 1361 -105
rect 1327 -313 1361 -297
rect 1423 -121 1457 -105
rect 1423 -313 1457 -297
rect 1519 -121 1553 -105
rect 1519 -313 1553 -297
rect 1615 -121 1649 -105
rect 1615 -313 1649 -297
rect 1711 -121 1745 -105
rect 1711 -313 1745 -297
rect 1807 -121 1841 -105
rect 1807 -313 1841 -297
rect 1903 -121 1937 -105
rect 1903 -313 1937 -297
rect 2017 -449 2051 -387
rect -2051 -483 -1955 -449
rect 1955 -483 2051 -449
<< viali >>
rect -1937 121 -1903 297
rect -1841 121 -1807 297
rect -1745 121 -1711 297
rect -1649 121 -1615 297
rect -1553 121 -1519 297
rect -1457 121 -1423 297
rect -1361 121 -1327 297
rect -1265 121 -1231 297
rect -1169 121 -1135 297
rect -1073 121 -1039 297
rect -977 121 -943 297
rect -881 121 -847 297
rect -785 121 -751 297
rect -689 121 -655 297
rect -593 121 -559 297
rect -497 121 -463 297
rect -401 121 -367 297
rect -305 121 -271 297
rect -209 121 -175 297
rect -113 121 -79 297
rect -17 121 17 297
rect 79 121 113 297
rect 175 121 209 297
rect 271 121 305 297
rect 367 121 401 297
rect 463 121 497 297
rect 559 121 593 297
rect 655 121 689 297
rect 751 121 785 297
rect 847 121 881 297
rect 943 121 977 297
rect 1039 121 1073 297
rect 1135 121 1169 297
rect 1231 121 1265 297
rect 1327 121 1361 297
rect 1423 121 1457 297
rect 1519 121 1553 297
rect 1615 121 1649 297
rect 1711 121 1745 297
rect 1807 121 1841 297
rect 1903 121 1937 297
rect -1937 -297 -1903 -121
rect -1841 -297 -1807 -121
rect -1745 -297 -1711 -121
rect -1649 -297 -1615 -121
rect -1553 -297 -1519 -121
rect -1457 -297 -1423 -121
rect -1361 -297 -1327 -121
rect -1265 -297 -1231 -121
rect -1169 -297 -1135 -121
rect -1073 -297 -1039 -121
rect -977 -297 -943 -121
rect -881 -297 -847 -121
rect -785 -297 -751 -121
rect -689 -297 -655 -121
rect -593 -297 -559 -121
rect -497 -297 -463 -121
rect -401 -297 -367 -121
rect -305 -297 -271 -121
rect -209 -297 -175 -121
rect -113 -297 -79 -121
rect -17 -297 17 -121
rect 79 -297 113 -121
rect 175 -297 209 -121
rect 271 -297 305 -121
rect 367 -297 401 -121
rect 463 -297 497 -121
rect 559 -297 593 -121
rect 655 -297 689 -121
rect 751 -297 785 -121
rect 847 -297 881 -121
rect 943 -297 977 -121
rect 1039 -297 1073 -121
rect 1135 -297 1169 -121
rect 1231 -297 1265 -121
rect 1327 -297 1361 -121
rect 1423 -297 1457 -121
rect 1519 -297 1553 -121
rect 1615 -297 1649 -121
rect 1711 -297 1745 -121
rect 1807 -297 1841 -121
rect 1903 -297 1937 -121
<< metal1 >>
rect -1943 297 -1897 309
rect -1943 121 -1937 297
rect -1903 121 -1897 297
rect -1943 109 -1897 121
rect -1847 297 -1801 309
rect -1847 121 -1841 297
rect -1807 121 -1801 297
rect -1847 109 -1801 121
rect -1751 297 -1705 309
rect -1751 121 -1745 297
rect -1711 121 -1705 297
rect -1751 109 -1705 121
rect -1655 297 -1609 309
rect -1655 121 -1649 297
rect -1615 121 -1609 297
rect -1655 109 -1609 121
rect -1559 297 -1513 309
rect -1559 121 -1553 297
rect -1519 121 -1513 297
rect -1559 109 -1513 121
rect -1463 297 -1417 309
rect -1463 121 -1457 297
rect -1423 121 -1417 297
rect -1463 109 -1417 121
rect -1367 297 -1321 309
rect -1367 121 -1361 297
rect -1327 121 -1321 297
rect -1367 109 -1321 121
rect -1271 297 -1225 309
rect -1271 121 -1265 297
rect -1231 121 -1225 297
rect -1271 109 -1225 121
rect -1175 297 -1129 309
rect -1175 121 -1169 297
rect -1135 121 -1129 297
rect -1175 109 -1129 121
rect -1079 297 -1033 309
rect -1079 121 -1073 297
rect -1039 121 -1033 297
rect -1079 109 -1033 121
rect -983 297 -937 309
rect -983 121 -977 297
rect -943 121 -937 297
rect -983 109 -937 121
rect -887 297 -841 309
rect -887 121 -881 297
rect -847 121 -841 297
rect -887 109 -841 121
rect -791 297 -745 309
rect -791 121 -785 297
rect -751 121 -745 297
rect -791 109 -745 121
rect -695 297 -649 309
rect -695 121 -689 297
rect -655 121 -649 297
rect -695 109 -649 121
rect -599 297 -553 309
rect -599 121 -593 297
rect -559 121 -553 297
rect -599 109 -553 121
rect -503 297 -457 309
rect -503 121 -497 297
rect -463 121 -457 297
rect -503 109 -457 121
rect -407 297 -361 309
rect -407 121 -401 297
rect -367 121 -361 297
rect -407 109 -361 121
rect -311 297 -265 309
rect -311 121 -305 297
rect -271 121 -265 297
rect -311 109 -265 121
rect -215 297 -169 309
rect -215 121 -209 297
rect -175 121 -169 297
rect -215 109 -169 121
rect -119 297 -73 309
rect -119 121 -113 297
rect -79 121 -73 297
rect -119 109 -73 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 73 297 119 309
rect 73 121 79 297
rect 113 121 119 297
rect 73 109 119 121
rect 169 297 215 309
rect 169 121 175 297
rect 209 121 215 297
rect 169 109 215 121
rect 265 297 311 309
rect 265 121 271 297
rect 305 121 311 297
rect 265 109 311 121
rect 361 297 407 309
rect 361 121 367 297
rect 401 121 407 297
rect 361 109 407 121
rect 457 297 503 309
rect 457 121 463 297
rect 497 121 503 297
rect 457 109 503 121
rect 553 297 599 309
rect 553 121 559 297
rect 593 121 599 297
rect 553 109 599 121
rect 649 297 695 309
rect 649 121 655 297
rect 689 121 695 297
rect 649 109 695 121
rect 745 297 791 309
rect 745 121 751 297
rect 785 121 791 297
rect 745 109 791 121
rect 841 297 887 309
rect 841 121 847 297
rect 881 121 887 297
rect 841 109 887 121
rect 937 297 983 309
rect 937 121 943 297
rect 977 121 983 297
rect 937 109 983 121
rect 1033 297 1079 309
rect 1033 121 1039 297
rect 1073 121 1079 297
rect 1033 109 1079 121
rect 1129 297 1175 309
rect 1129 121 1135 297
rect 1169 121 1175 297
rect 1129 109 1175 121
rect 1225 297 1271 309
rect 1225 121 1231 297
rect 1265 121 1271 297
rect 1225 109 1271 121
rect 1321 297 1367 309
rect 1321 121 1327 297
rect 1361 121 1367 297
rect 1321 109 1367 121
rect 1417 297 1463 309
rect 1417 121 1423 297
rect 1457 121 1463 297
rect 1417 109 1463 121
rect 1513 297 1559 309
rect 1513 121 1519 297
rect 1553 121 1559 297
rect 1513 109 1559 121
rect 1609 297 1655 309
rect 1609 121 1615 297
rect 1649 121 1655 297
rect 1609 109 1655 121
rect 1705 297 1751 309
rect 1705 121 1711 297
rect 1745 121 1751 297
rect 1705 109 1751 121
rect 1801 297 1847 309
rect 1801 121 1807 297
rect 1841 121 1847 297
rect 1801 109 1847 121
rect 1897 297 1943 309
rect 1897 121 1903 297
rect 1937 121 1943 297
rect 1897 109 1943 121
rect -1943 -121 -1897 -109
rect -1943 -297 -1937 -121
rect -1903 -297 -1897 -121
rect -1943 -309 -1897 -297
rect -1847 -121 -1801 -109
rect -1847 -297 -1841 -121
rect -1807 -297 -1801 -121
rect -1847 -309 -1801 -297
rect -1751 -121 -1705 -109
rect -1751 -297 -1745 -121
rect -1711 -297 -1705 -121
rect -1751 -309 -1705 -297
rect -1655 -121 -1609 -109
rect -1655 -297 -1649 -121
rect -1615 -297 -1609 -121
rect -1655 -309 -1609 -297
rect -1559 -121 -1513 -109
rect -1559 -297 -1553 -121
rect -1519 -297 -1513 -121
rect -1559 -309 -1513 -297
rect -1463 -121 -1417 -109
rect -1463 -297 -1457 -121
rect -1423 -297 -1417 -121
rect -1463 -309 -1417 -297
rect -1367 -121 -1321 -109
rect -1367 -297 -1361 -121
rect -1327 -297 -1321 -121
rect -1367 -309 -1321 -297
rect -1271 -121 -1225 -109
rect -1271 -297 -1265 -121
rect -1231 -297 -1225 -121
rect -1271 -309 -1225 -297
rect -1175 -121 -1129 -109
rect -1175 -297 -1169 -121
rect -1135 -297 -1129 -121
rect -1175 -309 -1129 -297
rect -1079 -121 -1033 -109
rect -1079 -297 -1073 -121
rect -1039 -297 -1033 -121
rect -1079 -309 -1033 -297
rect -983 -121 -937 -109
rect -983 -297 -977 -121
rect -943 -297 -937 -121
rect -983 -309 -937 -297
rect -887 -121 -841 -109
rect -887 -297 -881 -121
rect -847 -297 -841 -121
rect -887 -309 -841 -297
rect -791 -121 -745 -109
rect -791 -297 -785 -121
rect -751 -297 -745 -121
rect -791 -309 -745 -297
rect -695 -121 -649 -109
rect -695 -297 -689 -121
rect -655 -297 -649 -121
rect -695 -309 -649 -297
rect -599 -121 -553 -109
rect -599 -297 -593 -121
rect -559 -297 -553 -121
rect -599 -309 -553 -297
rect -503 -121 -457 -109
rect -503 -297 -497 -121
rect -463 -297 -457 -121
rect -503 -309 -457 -297
rect -407 -121 -361 -109
rect -407 -297 -401 -121
rect -367 -297 -361 -121
rect -407 -309 -361 -297
rect -311 -121 -265 -109
rect -311 -297 -305 -121
rect -271 -297 -265 -121
rect -311 -309 -265 -297
rect -215 -121 -169 -109
rect -215 -297 -209 -121
rect -175 -297 -169 -121
rect -215 -309 -169 -297
rect -119 -121 -73 -109
rect -119 -297 -113 -121
rect -79 -297 -73 -121
rect -119 -309 -73 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 73 -121 119 -109
rect 73 -297 79 -121
rect 113 -297 119 -121
rect 73 -309 119 -297
rect 169 -121 215 -109
rect 169 -297 175 -121
rect 209 -297 215 -121
rect 169 -309 215 -297
rect 265 -121 311 -109
rect 265 -297 271 -121
rect 305 -297 311 -121
rect 265 -309 311 -297
rect 361 -121 407 -109
rect 361 -297 367 -121
rect 401 -297 407 -121
rect 361 -309 407 -297
rect 457 -121 503 -109
rect 457 -297 463 -121
rect 497 -297 503 -121
rect 457 -309 503 -297
rect 553 -121 599 -109
rect 553 -297 559 -121
rect 593 -297 599 -121
rect 553 -309 599 -297
rect 649 -121 695 -109
rect 649 -297 655 -121
rect 689 -297 695 -121
rect 649 -309 695 -297
rect 745 -121 791 -109
rect 745 -297 751 -121
rect 785 -297 791 -121
rect 745 -309 791 -297
rect 841 -121 887 -109
rect 841 -297 847 -121
rect 881 -297 887 -121
rect 841 -309 887 -297
rect 937 -121 983 -109
rect 937 -297 943 -121
rect 977 -297 983 -121
rect 937 -309 983 -297
rect 1033 -121 1079 -109
rect 1033 -297 1039 -121
rect 1073 -297 1079 -121
rect 1033 -309 1079 -297
rect 1129 -121 1175 -109
rect 1129 -297 1135 -121
rect 1169 -297 1175 -121
rect 1129 -309 1175 -297
rect 1225 -121 1271 -109
rect 1225 -297 1231 -121
rect 1265 -297 1271 -121
rect 1225 -309 1271 -297
rect 1321 -121 1367 -109
rect 1321 -297 1327 -121
rect 1361 -297 1367 -121
rect 1321 -309 1367 -297
rect 1417 -121 1463 -109
rect 1417 -297 1423 -121
rect 1457 -297 1463 -121
rect 1417 -309 1463 -297
rect 1513 -121 1559 -109
rect 1513 -297 1519 -121
rect 1553 -297 1559 -121
rect 1513 -309 1559 -297
rect 1609 -121 1655 -109
rect 1609 -297 1615 -121
rect 1649 -297 1655 -121
rect 1609 -309 1655 -297
rect 1705 -121 1751 -109
rect 1705 -297 1711 -121
rect 1745 -297 1751 -121
rect 1705 -309 1751 -297
rect 1801 -121 1847 -109
rect 1801 -297 1807 -121
rect 1841 -297 1847 -121
rect 1801 -309 1847 -297
rect 1897 -121 1943 -109
rect 1897 -297 1903 -121
rect 1937 -297 1943 -121
rect 1897 -309 1943 -297
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -2034 -466 2034 466
string parameters w 1 l 0.150 m 2 nf 40 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
