magic
tech sky130A
magscale 1 2
timestamp 1623980668
<< pwell >>
rect -226 -321 226 510
rect -226 -387 -114 -321
rect -48 -322 226 -321
rect -226 -388 -111 -387
rect -99 -388 226 -322
rect -226 -510 226 -388
<< nmos >>
rect -30 -300 30 300
<< ndiff >>
rect -88 288 -30 300
rect -88 -288 -76 288
rect -42 -288 -30 288
rect -88 -300 -30 -288
rect 30 288 88 300
rect 30 -288 42 288
rect 76 -288 88 288
rect 30 -300 88 -288
<< ndiffc >>
rect -76 -288 -42 288
rect 42 -288 76 288
<< psubdiff >>
rect -190 440 -94 474
rect 94 440 190 474
rect -190 378 -156 440
rect 156 378 190 440
rect -190 -440 -156 -378
rect 156 -440 190 -378
rect -190 -474 -94 -440
rect 94 -474 190 -440
<< psubdiffcont >>
rect -94 440 94 474
rect -190 -378 -156 378
rect 156 -378 190 378
rect -94 -474 94 -440
<< poly >>
rect -30 300 30 326
rect -30 -322 30 -300
rect -99 -338 33 -322
rect -99 -372 -83 -338
rect 17 -372 33 -338
rect -99 -388 33 -372
<< polycont >>
rect -83 -372 17 -338
<< locali >>
rect -190 440 -94 474
rect 94 440 190 474
rect -190 378 -156 440
rect 156 378 190 440
rect -76 288 -42 304
rect -76 -304 -42 -288
rect 42 288 76 304
rect 42 -304 76 -288
rect -99 -372 -83 -338
rect 17 -372 33 -338
rect -190 -440 -156 -378
rect 156 -440 190 -378
rect -190 -474 -94 -440
rect 94 -474 190 -440
<< viali >>
rect -76 -288 -42 288
rect 42 -288 76 288
rect -83 -372 17 -338
<< metal1 >>
rect -82 288 -36 300
rect -82 -288 -76 288
rect -42 -288 -36 288
rect -82 -300 -36 -288
rect 36 288 82 300
rect 36 -288 42 288
rect 76 -288 82 288
rect 36 -300 82 -288
rect -98 -338 32 -329
rect -98 -372 -83 -338
rect 17 -372 32 -338
rect -98 -381 32 -372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -173 -457 173 457
string parameters w 3 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
